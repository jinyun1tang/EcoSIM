netcdf ecosim_pftpar_20251018 {
dimensions:
	npfts = UNLIMITED ; // (76 currently)
	JLI = 4 ;
	nchars1 = 10 ;
	npft = 35 ;
	nchars2 = 4 ;
	nchars3 = 40 ;
	nkopenclms = 31 ;
	nchars4 = 2 ;
	nchars5 = 3 ;
	nchars6 = 64 ;
variables:
	byte ICTYP(npfts) ;
		ICTYP:long_name = "photosynthesis type" ;
		ICTYP:units = "none" ;
		ICTYP:flags = "C3 or C4" ;
	byte IGTYP(npfts) ;
		IGTYP:long_name = "root profile" ;
		IGTYP:units = "none" ;
		IGTYP:flags = "0=shallow (eg bryophytes),1=intermediate(eg herbs),2=deep (eg trees)" ;
	byte ISTYP(npfts) ;
		ISTYP:long_name = "growth habit" ;
		ISTYP:units = "none" ;
		ISTYP:flags = "0=annual,1=perennial" ;
	byte IDTYP(npfts) ;
		IDTYP:long_name = "growth pattern" ;
		IDTYP:units = "none" ;
		IDTYP:flags = "0=determinate,1=indetermimate" ;
	byte INTYP(npfts) ;
		INTYP:long_name = "N2 fixation" ;
		INTYP:units = "none" ;
		INTYP:flags = "1,2,3=rapid to slow root symbiosis (e.g.legumes),4,5,6=rapid to slow canopy symbiosis (e.g. cyanobacteria)" ;
	byte IWTYP(npfts) ;
		IWTYP:long_name = "phenology type" ;
		IWTYP:units = "none" ;
		IWTYP:flags = "0=evergreen,1=cold deciduous,2=drought deciduous,3=1+2" ;
	byte IPTYP(npfts) ;
		IPTYP:long_name = "photoperiod type" ;
		IPTYP:units = "none" ;
		IPTYP:flags = "0=day neutral,1=short day,2=long day" ;
	byte IBTYP(npfts) ;
		IBTYP:long_name = "turnover of aboveground biomass" ;
		IBTYP:units = "none" ;
		IBTYP:flags = "0,1=rapid(fully deciduous),2=very slow(needle evergreen),3=(broadleaf evergreen),4=slow(semi-deciduous),5=(semi-evergreen)" ;
	byte IRTYP(npfts) ;
		IRTYP:long_name = "storage organ" ;
		IRTYP:units = "none" ;
		IRTYP:flags = "0=above ground,1=below ground" ;
	byte MY(npfts) ;
		MY:long_name = "mycorrhizal" ;
		MY:units = "none" ;
		MY:flags = "1=no,2=yes" ;
	float ZTYPI(npfts) ;
		ZTYPI:long_name = "thermal adaptation zone" ;
		ZTYPI:units = "none" ;
		ZTYPI:flags = "1=arctic,boreal,2=cool temperate" ;
	float VCMX(npfts) ;
		VCMX:long_name = "specific C3 rubisco carboxylase" ;
		VCMX:units = "umol C g-1 s-1" ;
	float VOMX(npfts) ;
		VOMX:long_name = "specific rubisco oxygenase activity" ;
		VOMX:units = "umol O g-1 s-1" ;
	float VCMX4(npfts) ;
		VCMX4:long_name = "specific PEP carboxylase activity" ;
		VCMX4:units = "umol g-1 s-1" ;
	float XKCO2(npfts) ;
		XKCO2:long_name = "Km for VCMX" ;
		XKCO2:units = "uM" ;
	float XKO2(npfts) ;
		XKO2:long_name = "Km for VOMX" ;
		XKO2:units = "uM" ;
	float XKCO24(npfts) ;
		XKCO24:long_name = "Km for VCMX4" ;
		XKCO24:units = "uM" ;
	float RUBP(npfts) ;
		RUBP:long_name = "fraction of leaf protein in rubisco" ;
		RUBP:units = "none" ;
	float PEPC(npfts) ;
		PEPC:long_name = "fraction of leaf protein in PEP carboxylase" ;
		PEPC:units = "none" ;
	float ETMX(npfts) ;
		ETMX:long_name = "specific chlorophyll activity" ;
		ETMX:units = "umol e- g-1 s-1" ;
	float CHL(npfts) ;
		CHL:long_name = "fraction of leaf protein in mesophyll(C3) chlorophyll" ;
		CHL:units = "none" ;
	float CHL4(npfts) ;
		CHL4:long_name = "fraction of leaf protein in bundle sheath(C4) chlorophyll" ;
		CHL4:units = "none" ;
	float FCO2(npfts) ;
		FCO2:long_name = "intercellular" ;
		FCO2:units = "none" ;
		FCO2:flags = "atmospheric CO2 concentration ratio" ;
	float ALBR(npfts) ;
		ALBR:long_name = "leaf SW albedo" ;
		ALBR:units = "none" ;
	float ALBP(npfts) ;
		ALBP:long_name = "leaf PAR albedo" ;
		ALBP:units = "none" ;
	float TAUR(npfts) ;
		TAUR:long_name = "leaf SW transmission" ;
		TAUR:units = "none" ;
	float TAUP(npfts) ;
		TAUP:long_name = "leaf PAR transmission" ;
		TAUP:units = "none" ;
	float XRNI(npfts) ;
		XRNI:long_name = "rate of node initiation at 25oC" ;
		XRNI:units = "h-1" ;
	float XRLA(npfts) ;
		XRLA:long_name = "rate of leaf appearance at 25oC" ;
		XRLA:units = "h-1" ;
	float CTC(npfts) ;
		CTC:long_name = "chilling temperature for CO2 fixation, seed loss" ;
		CTC:units = "oC" ;
	float VRNLI(npfts) ;
		VRNLI:long_name = "hour requirement for spring leafout" ;
		VRNLI:units = "h" ;
	float VRNXI(npfts) ;
		VRNXI:long_name = "hour requirement for autumn leafoff" ;
		VRNXI:units = "h" ;
	float WDLF(npfts) ;
		WDLF:long_name = "leaf length vs width ratio" ;
		WDLF:units = "none" ;
	float PB(npfts) ;
		PB:long_name = "nonstructural C concentration needed for branching" ;
		PB:units = "gC gC-1" ;
	float GROUPX(npfts) ;
		GROUPX:long_name = "initial plant maturity group, aka minimum number of vegetative nodes initiated before floral" ;
		GROUPX:units = "none" ;
	float XTLI(npfts) ;
		XTLI:long_name = "node number in seed at planting" ;
		XTLI:units = "none" ;
	float XDL(npfts) ;
		XDL:long_name = "critical daylength for phenological progress" ;
		XDL:units = "h" ;
	float XPPD(npfts) ;
		XPPD:long_name = "photoperiod sensitivity, i.e. difference between current and critical daylengths used to calculate  phenological progress" ;
		XPPD:units = "node h-1" ;
	float SLA1(npfts) ;
		SLA1:long_name = "growth in leaf area vs mass" ;
		SLA1:units = "m2 gC-1" ;
	float SSL1(npfts) ;
		SSL1:long_name = "growth in petiole length vs mass" ;
		SSL1:units = "m gC-1" ;
	float SNL1(npfts) ;
		SNL1:long_name = "growth in internode stalk length vs mass" ;
		SNL1:units = "m gC-1" ;
	float CLASS(npfts, JLI) ;
		CLASS:long_name = "fraction of leaf area in 0-22.5,45,67.5,90o inclination classes" ;
		CLASS:units = "none" ;
	float CFI(npfts) ;
		CFI:long_name = "initial clumping factor" ;
		CFI:units = "none" ;
	float ANGBR(npfts) ;
		ANGBR:long_name = "stem angle from horizontal" ;
		ANGBR:units = "degree" ;
	float ANGSH(npfts) ;
		ANGSH:long_name = "petiole angle from horizontal" ;
		ANGSH:units = "degree" ;
	float STMX(npfts) ;
		STMX:long_name = "maximum potential seed sites for pre-anthesis stalk growth" ;
		STMX:units = "sites gC-1" ;
	float SDMX(npfts) ;
		SDMX:long_name = "maximum seed number per site" ;
		SDMX:units = "seeds site-1" ;
	float GRMX(npfts) ;
		GRMX:long_name = "maximum seed size per seed" ;
		GRMX:units = "gC seed-1" ;
	float GRDM(npfts) ;
		GRDM:long_name = "seed size at planting" ;
		GRDM:units = "gC seed-1" ;
	float GFILL(npfts) ;
		GFILL:long_name = "grain filling rate at 25 oC" ;
		GFILL:units = "gC seed-1 h-1" ;
	float WTSTDI(npfts) ;
		WTSTDI:long_name = "mass of dead standing biomass at planting" ;
		WTSTDI:units = "gC m-2" ;
	float RRAD1M(npfts) ;
		RRAD1M:long_name = "radius of primary root tips" ;
		RRAD1M:units = "m" ;
	float RRAD2M(npfts) ;
		RRAD2M:long_name = "radius of secondary roots" ;
		RRAD2M:units = "m" ;
	float PORT(npfts) ;
		PORT:long_name = "root porosity" ;
		PORT:units = "m3 m-3" ;
	float PR(npfts) ;
		PR:long_name = "nonstructural C concentration needed for root branching" ;
		PR:units = "gC gC-1" ;
	float RSRR(npfts) ;
		RSRR:long_name = "radial root resistivity" ;
		RSRR:units = "m2 MPa-1 h-1" ;
	float RSRA(npfts) ;
		RSRA:long_name = "axial root resistivity" ;
		RSRA:units = "m2 MPa-1 h-1" ;
	float PTSHT(npfts) ;
		PTSHT:long_name = "rate constant for equilibrating shoot-root nonstructural C concentration" ;
		PTSHT:units = "h-1" ;
	float RTFQ(npfts) ;
		RTFQ:long_name = "root branching frequency" ;
		RTFQ:units = "m-1" ;
	float UPMXZH(npfts) ;
		UPMXZH:long_name = "NH4 max uptake" ;
		UPMXZH:units = "g m-2 h-1" ;
	float UPKMZH(npfts) ;
		UPKMZH:long_name = "NH4 uptake Km" ;
		UPKMZH:units = "uM" ;
	float UPMNZH(npfts) ;
		UPMNZH:long_name = "NH4 uptake minimum conconcentration" ;
		UPMNZH:units = "uM" ;
	float UPMXZO(npfts) ;
		UPMXZO:long_name = "NO3 max uptake" ;
		UPMXZO:units = "g m-2 h-1" ;
	float UPKMZO(npfts) ;
		UPKMZO:long_name = "NO3 uptake Km" ;
		UPKMZO:units = "uM" ;
	float UPMNZO(npfts) ;
		UPMNZO:long_name = "NO3 uptake minimum conconcentration" ;
		UPMNZO:units = "uM" ;
	float UPMXPO(npfts) ;
		UPMXPO:long_name = "H2PO4 max uptake" ;
		UPMXPO:units = "gP m-2 h-1" ;
	float UPKMPO(npfts) ;
		UPKMPO:long_name = "H2PO4 uptake Km" ;
		UPKMPO:units = "uM" ;
	float UPMNPO(npfts) ;
		UPMNPO:long_name = "H2PO4 uptake minimum conconcentration" ;
		UPMNPO:units = "uM" ;
	float OSMO(npfts) ;
		OSMO:long_name = "leaf osmotic potential at zero leaf water potential" ;
		OSMO:units = "MPa" ;
	float RCS(npfts) ;
		RCS:long_name = "e-folding turgor pressure for stomatal resistance" ;
		RCS:units = "MPa" ;
	float RSMX(npfts) ;
		RSMX:long_name = "cuticular resistance" ;
		RSMX:units = "s m-1" ;
	float DMLF(npfts) ;
		DMLF:long_name = "leaf dry matter C production vs nonstructural C consumption" ;
		DMLF:units = "gC gC-1" ;
	float DMSHE(npfts) ;
		DMSHE:long_name = "petiole dry matter C production vs nonstructural C consumption" ;
		DMSHE:units = "gC gC-1" ;
	float DMSTK(npfts) ;
		DMSTK:long_name = "stalk dry matter C production vs nonstructural C consumption" ;
		DMSTK:units = "gC gC-1" ;
	float DMRSV(npfts) ;
		DMRSV:long_name = "stalk reserve C production vs nonstructural C consumption" ;
		DMRSV:units = "gC gC-1)" ;
	float DMHSK(npfts) ;
		DMHSK:long_name = "husk dry matter C production vs nonstructural Cconsumption" ;
		DMHSK:units = "gC gC-1" ;
	float DMEAR(npfts) ;
		DMEAR:long_name = "ear dry matter C production vs nonstructural Cconsumption" ;
		DMEAR:units = "gC gC-1" ;
	float DMGR(npfts) ;
		DMGR:long_name = "grain C production vs nonstructural C consumption" ;
		DMGR:units = "gC gC-1" ;
	float DMRT(npfts) ;
		DMRT:long_name = "root dry matter C production vs nonstructural C consumption" ;
		DMRT:units = "gC gC-1" ;
	float DMND(npfts) ;
		DMND:long_name = "nodule bacteria in root nodule,canopy dry matter C production vs nonstructural C consumption" ;
		DMND:units = "gC gC-1" ;
	float CNWR(npfts) ;
		CNWR:long_name = "Protein C to root N ratio in plant roots" ;
		CNWR:units = "gC gN-1" ;
	float CNWL(npfts) ;
		CNWL:long_name = "Protein C to leaf N ratio in plant leaves" ;
		CNWL:units = "gC gN-1" ;
	float CNLF(npfts) ;
		CNLF:long_name = "NC ratio in plant leaves" ;
		CNLF:units = "gN gC-1" ;
	float CNSHE(npfts) ;
		CNSHE:long_name = "NC ratio in plant petiole" ;
		CNSHE:units = "gN gC-1" ;
	float CNSTK(npfts) ;
		CNSTK:long_name = "NC ratio in plant stalk" ;
		CNSTK:units = "gN gC-1" ;
	float CNRSV(npfts) ;
		CNRSV:long_name = "NC ratio in plant stalk reserve" ;
		CNRSV:units = "gN gC-1" ;
	float CNHSK(npfts) ;
		CNHSK:long_name = "NC ratio in plant husk" ;
		CNHSK:units = "gN gC-1" ;
	float CNEAR(npfts) ;
		CNEAR:long_name = "NC ratio in plant ear" ;
		CNEAR:units = "gN gC-1" ;
	float CNGR(npfts) ;
		CNGR:long_name = "NC ratio in plant grain" ;
		CNGR:units = "gN gC-1" ;
	float CNRT(npfts) ;
		CNRT:long_name = "NC ratio in plant root" ;
		CNRT:units = "gN gC-1" ;
	float CNND(npfts) ;
		CNND:long_name = "NC ratio in plant nodule" ;
		CNND:units = "gN gC-1" ;
	float CPWR(npfts) ;
		CPWR:long_name = "Protein C to root P ratio in plant roots" ;
		CPWR:units = "gC gP-1" ;
	float CPWL(npfts) ;
		CPWL:long_name = "Protein C to leaf P ratio in plant leaves" ;
		CPWL:units = "gC gP-1" ;
	float CPLF(npfts) ;
		CPLF:long_name = "PC ratio in plant leaves" ;
		CPLF:units = "gP gC-1" ;
	float CPSHE(npfts) ;
		CPSHE:long_name = "PC ratio in plant petiole" ;
		CPSHE:units = "gP gC-1" ;
	float CPSTK(npfts) ;
		CPSTK:long_name = "PC ratio in plant stalk" ;
		CPSTK:units = "gP gC-1" ;
	float CPRSV(npfts) ;
		CPRSV:long_name = "PC ratio in plant stalk reserve" ;
		CPRSV:units = "gP gC-1" ;
	float CPHSK(npfts) ;
		CPHSK:long_name = "PC ratio in plant husk" ;
		CPHSK:units = "gP gC-1" ;
	float CPEAR(npfts) ;
		CPEAR:long_name = "PC ratio in plant ear" ;
		CPEAR:units = "gP gC-1" ;
	float CPGR(npfts) ;
		CPGR:long_name = "PC ratio in plant grain" ;
		CPGR:units = "gP gC-1" ;
	float CPRT(npfts) ;
		CPRT:long_name = "PC ratio in plant root" ;
		CPRT:units = "gP gC-1" ;
	float CPND(npfts) ;
		CPND:long_name = "PC ratio in plant nodule" ;
		CPND:units = "gP gC-1" ;
   float ROOTMAGE(npfts) ;
      ROOTMAGE:long_name="Root maturation age to trigger secondary growth" ;
      ROOTMAGE:units ="h" ;
	char pfts(npfts, nchars1) ;
	char pfts_short(npft, nchars2) ;
	char pfts_long(npft, nchars3) ;
	char koppen_clim_no(nkopenclms, nchars4) ;
	char koppen_clim_short(nkopenclms, nchars5) ;
	char koppen_clim_long(nkopenclms, nchars6) ;

// global attributes:
		:description = "plant trait parameterization for ecosim created on 2024/03/14/10:02:16" ;
		:history = "Sat Oct 18 12:06:29 2025: ncrcat ecosim_pftpar_20240723.nc /Users/jinyuntang/work/github/ecosim_benchmark/RiceUSTWT/Rice_pftpar_20251017.nc ecosim_pftpar_20251018.nc" ;
		:NCO = "netCDF Operators version 5.3.5 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 ICTYP = 3, 3, 3, 3, 4, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 
    3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 4, 3, 3, 3, 3, 
    3, 3, 4, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 
    3, 3, 3, 3, 3 ;

 IGTYP = 1, 1, 2, 1, 1, 0, 3, 1, 2, 1, 0, 3, 1, 1, 1, 0, 2, 1, 2, 2, 2, 2, 2, 
    1, 2, 2, 2, 2, 3, 1, 2, 2, 3, 3, 1, 2, 1, 0, 1, 0, 1, 1, 1, 1, 0, 2, 0, 
    2, 2, 1, 3, 2, 2, 1, 2, 1, 2, 2, 1, 2, 1, 3, 2, 2, 0, 1, 3, 0, 1, 0, 0, 
    0, 1, 3, 1, 1 ;

 ISTYP = 1, 1, 1, 1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 1, 0, 0, 1, 1, 
    0, 1, 1, 1, 1, 1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0, 1, 1, 1, 0, 0, 1, 1, 1, 0, 1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0, 1, 0, 0 ;

 IDTYP = 0, 0, 1, 0, 0, 1, 1, 0, 1, 0, 1, 1, 0, 1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0, 1, 1, 1, 1, 1, 1, 0, 1, 0, 1, 0, 1, 0, 0, 1, 1, 1, 
    1, 1, 0, 1, 1, 1, 0, 1, 1, 1, 1, 0, 1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0, 1, 1, 0 ;

 INTYP = 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 4, 1, 0, 2, 1, 6, 0, 0, 0, 1, 2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 2, 0, 0, 5, 0, 5, 0, 0, 0, 0, 5, 2, 6, 
    0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 2, 0, 0, 0, 0, 0, 3, 3, 3, 0, 3, 2, 5, 5, 
    6, 0, 0, 0, 0 ;

 IWTYP = 1, 1, 1, 1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 2, 0, 0, 2, 1, 1, 
    2, 1, 0, 0, 1, 1, 0, 1, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0, 0, 0, 1, 1, 0, 0, 1, 1, 1, 0, 1, 0, 0, 1, 0, 1, 1, 1, 1, 1, 1, 1, 
    1, 0, 0, 2, 0 ;

 IPTYP = 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 2, 2, 2, 2, 2, 2, 
    2, 2, 0, 0, 2, 2, 0, 2, 2, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 2, 0, 2, 2, 0, 2, 2, 2, 2, 2, 2, 0, 
    2, 1, 2, 2, 0 ;

 IBTYP = 0, 0, 0, 0, 0, 2, 2, 0, 0, 0, 2, 0, 0, 0, 0, 3, 3, 0, 2, 0, 0, 1, 1, 
    0, 1, 2, 2, 1, 2, 0, 1, 2, 2, 0, 0, 2, 0, 3, 0, 3, 0, 0, 0, 0, 3, 0, 3, 
    2, 2, 0, 2, 1, 1, 0, 0, 0, 1, 1, 0, 1, 0, 2, 2, 1, 2, 0, 1, 2, 0, 3, 3, 
    3, 0, 2, 0, 0 ;

 IRTYP = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0 ;

 MY = 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2 ;

 ZTYPI = 1, 1.5, 3, 1, 2.5, 1, 1, 1, 2.5, 1, 1, 1, 1, 1.5, 1.5, 1, 5, 2, 1, 
    2.5, 2, 1, 1, 2, 1, 1.5, 3, 1.5, 1, 2, 2, 3, 1.5, 1.5, 1, 1, 1, 1, 1.5, 
    1, 1.2, 1.5, 1.5, 1, 1, 3, 1, 1, 1.5, 1.5, 3, 1, 1, 1.5, 1.5, 1, 3, 1.5, 
    2, 1, 2, 3, 1, 5, 1, 1.5, 3, 1, 1, 1, 1, 1, 3, 3, 2, 2 ;

 VCMX = 45, 45, 45, 45, 60, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 
    30, 45, 50, 30, 45, 45, 45, 45, 45, 30, 45, 45, 45, 45, 45, 45, 45, 45, 
    45, 90, 45, 45, 45, 45, 45, 75, 45, 45, 45, 45, 45, 45, 90, 45, 45, 45, 
    45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 
    45, 250, 30, 25, 45 ;

 VOMX = 9.5, 9.5, 9.5, 9.5, 12, 9.5, 9.5, 9.5, 9.5, 9.5, 9.5, 9.5, 9.5, 9.5, 
    9.5, 9.5, 9.5, 9.5, 9.5, 12, 9.5, 9.5, 9.5, 9.5, 9.5, 9.5, 9.5, 9.5, 9.5, 
    9.5, 9.5, 9.5, 9.5, 9.5, 9.5, 9.5, 9.5, 9.5, 9.5, 9.5, 9.5, 9.5, 15, 9.5, 
    9.5, 9.5, 9.5, 9.5, 9.5, 15, 9.5, 9.5, 9.5, 9.5, 9.5, 9.5, 9.5, 9.5, 9.5, 
    9.5, 9.5, 9.5, 9.5, 9.5, 9.5, 9.5, 9.5, 9.5, 9.5, 9.5, 9.5, 9.5, 0.25, 
    9.5, 9.5, 9.5 ;

 VCMX4 = 0, 0, 0, 0, 900, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 150, 0, 0, 0, 
    0, 0, 0, 180, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0 ;

 XKCO2 = 12.5, 12.5, 12.5, 12.5, 30, 12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 
    12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 
    12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 
    12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 30, 12.5, 12.5, 12.5, 12.5, 
    12.5, 12.5, 30, 12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 
    12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 12.5, 
    12.5, 12.5, 12.5, 12.5, 12.5 ;

 XKO2 = 500, 500, 500, 500, 810, 500, 500, 500, 500, 500, 500, 500, 500, 500, 
    500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 
    500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 
    810, 500, 500, 500, 500, 500, 500, 810, 500, 500, 500, 500, 500, 500, 
    500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 
    500, 500, 400, 500, 500, 500 ;

 XKCO24 = 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0 ;

 RUBP = 0.125, 0.125, 0.125, 0.125, 0.1, 0.125, 0.125, 0.125, 0.125, 0.2, 
    0.125, 0.2, 0.125, 0.125, 0.125, 0.125, 0.125, 0.25, 0.125, 0.25, 0.25, 
    0.125, 0.125, 0.125, 0.125, 0.125, 0.125, 0.125, 0.125, 0.2, 0.125, 
    0.125, 0.125, 0.125, 0.125, 0.125, 0.125, 0.125, 0.125, 0.125, 0.125, 
    0.125, 0.025, 0.125, 0.125, 0.125, 0.125, 0.125, 0.125, 0.025, 0.125, 
    0.125, 0.125, 0.167, 0.167, 0.125, 0.125, 0.125, 0.2, 0.125, 0.2, 0.125, 
    0.125, 0.125, 0.125, 0.125, 0.125, 0.125, 0.125, 0.125, 0.125, 0.125, 
    0.3, 0.125, 0.25, 0.2 ;

 PEPC = 0, 0, 0, 0, 0.015, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.05, 0, 0, 
    0, 0, 0, 0, 0.05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0 ;

 ETMX = 405, 405, 405, 500, 600, 405, 405, 405, 450, 405, 405, 405, 405, 405, 
    405, 405, 405, 250, 405, 750, 250, 405, 405, 405, 405, 405, 320, 405, 
    405, 405, 405, 450, 405, 405, 405, 405, 500, 405, 405, 405, 405, 405, 
    405, 405, 405, 405, 405, 405, 405, 405, 405, 405, 405, 405, 405, 405, 
    405, 405, 405, 405, 405, 405, 405, 405, 405, 405, 405, 405, 405, 405, 
    405, 405, 500, 350, 220, 405 ;

 CHL = 0.025, 0.025, 0.025, 0.025, 0.1, 0.025, 0.025, 0.025, 0.025, 0.04, 
    0.025, 0.04, 0.025, 0.025, 0.025, 0.025, 0.025, 0.04, 0.025, 0.04, 0.04, 
    0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.04, 0.025, 
    0.025, 0.025, 0.025, 0.025, 0.025, 0.07, 0.025, 0.025, 0.025, 0.025, 
    0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 
    0.025, 0.025, 0.033, 0.033, 0.025, 0.025, 0.025, 0.04, 0.025, 0.04, 
    0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 0.025, 
    0.025, 0.04, 0.025, 0.04, 0.04 ;

 CHL4 = 0, 0, 0, 0, 0.15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.05, 0, 0, 
    0, 0, 0, 0, 0.05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0 ;

 FCO2 = 0.7, 0.7, 0.7, 0.8, 0.45, 0.7, 0.7, 0.7, 0.7, 0.7, 0.7, 0.7, 0.7, 
    0.7, 0.7, 0.7, 0.8, 0.7, 0.7, 0.7, 0.7, 0.7, 0.7, 0.7, 0.7, 0.7, 0.7, 
    0.7, 0.7, 0.7, 0.7, 0.75, 0.7, 0.7, 0.7, 0.7, 0.7, 0.7, 0.7, 0.7, 0.7, 
    0.7, 0.45, 0.7, 1, 0.7, 0.7, 0.7, 0.7, 0.45, 0.7, 0.7, 0.7, 0.7, 0.7, 
    0.7, 0.7, 0.7, 0.7, 0.7, 0.7, 0.7, 0.7, 0.75, 0.7, 0.7, 0.7, 0.7, 0.7, 
    0.7, 0.7, 1, 0.85, 0.7, 0.7, 0.7 ;

 ALBR = 0.15, 0.15, 0.15, 0.15, 0.2, 0.15, 0.15, 0.15, 0.15, 0.15, 0.15, 
    0.15, 0.15, 0.15, 0.15, 0.15, 0.15, 0.2, 0.09, 0.2, 0.2, 0.2, 0.15, 0.2, 
    0.15, 0.1, 0.125, 0.15, 0.1, 0.2, 0.15, 0.1, 0.1, 0.15, 0.15, 0.15, 0.15, 
    0.15, 0.15, 0.15, 0.15, 0.15, 0.15, 0.15, 0.2, 0.15, 0.15, 0.15, 0.15, 
    0.15, 0.15, 0.1, 0.15, 0.15, 0.15, 0.15, 0.15, 0.15, 0.2, 0.15, 0.2, 0.1, 
    0.15, 0.15, 0.15, 0.15, 0.15, 0.15, 0.15, 0.15, 0.15, 0.2, 0.2, 0.125, 
    0.2, 0.2 ;

 ALBP = 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.05, 0.075, 0.05, 0.075, 
    0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.05, 0.075, 0.05, 0.075, 
    0.075, 0.075, 0.075, 0.075, 0.075, 0.05, 0.05, 0.075, 0.05, 0.075, 0.075, 
    0.05, 0.05, 0.075, 0.075, 0.05, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 
    0.075, 0.075, 0.075, 0.075, 0.075, 0.05, 0.05, 0.075, 0.05, 0.05, 0.075, 
    0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.05, 0.075, 
    0.05, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 
    0.05, 0.075, 0.075 ;

 TAUR = 0.15, 0.15, 0.15, 0.15, 0.2, 0.15, 0.15, 0.15, 0.15, 0.15, 0.15, 
    0.15, 0.15, 0.15, 0.15, 0.15, 0.15, 0.2, 0.09, 0.2, 0.2, 0.2, 0.15, 0.2, 
    0.15, 0.1, 0.1, 0.15, 0.1, 0.2, 0.15, 0.1, 0.1, 0.15, 0.15, 0.15, 0.15, 
    0.15, 0.15, 0.15, 0.15, 0.15, 0.15, 0.15, 0.2, 0.15, 0.15, 0.15, 0.15, 
    0.15, 0.15, 0.1, 0.15, 0.15, 0.15, 0.15, 0.15, 0.15, 0.2, 0.15, 0.2, 0.1, 
    0.15, 0.15, 0.15, 0.15, 0.15, 0.15, 0.15, 0.15, 0.15, 0.2, 0.25, 0.15, 
    0.2, 0.2 ;

 TAUP = 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.05, 0.075, 0.05, 0.075, 
    0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.05, 0.075, 0.05, 0.075, 
    0.075, 0.075, 0.075, 0.075, 0.075, 0.05, 0.05, 0.075, 0.05, 0.075, 0.075, 
    0.05, 0.05, 0.075, 0.075, 0.05, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 
    0.075, 0.075, 0.075, 0.075, 0.075, 0.05, 0.05, 0.075, 0.05, 0.05, 0.075, 
    0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.05, 0.075, 
    0.05, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 
    0.05, 0.075, 0.075 ;

 XRNI = 0.015, 0.015, 0.015, 0.015, 0.025, 0.015, 0.015, 0.015, 0.015, 0.015, 
    0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.00225, 0.015, 
    0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 
    0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.00225, 0.015, 0.015, 0.015, 
    0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.025, 
    0.015, 0.015, 0.015, 0.015, 0.025, 0.015, 0.015, 0.015, 0.015, 0.015, 
    0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 0.015, 
    0.015, 0.015, 0.015, 0.015, 0.015, 0.015 ;

 XRLA = 0.009, 0.009, 0.009, 0.009, 0.015, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.0125, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.015, 
    0.009, 0.009, 0.009, 0.009, 0.015, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 0.009, 
    0.009, 0.009, 0.009, 0.009, 0.009, 0.009 ;

 CTC = -10, -5, 5, -10, 0, -10, -10, -20, 0, -10, -10, -10, -10, -5, -5, -20, 
    0, -5, -10, 0, -5, -10, -10, -5, -20, 0, 0, -5, -20, -10, -5, 0, 0, -5, 
    -10, -10, -10, -10, -5, -10, -10, -5, -5, -10, -10, 5, -10, -10, -7.5, 0, 
    0, -10, -10, -0.5, 0, -10, 0, 0, -10, -10, -10, 0, -10, 0, -10, -5, 0, 
    -10, -10, -10, -20, -10, 0, -7.5, -5, -5 ;

 VRNLI = 60, 360, 240, 40, 240, 60, 120, 48, 1500, 240, 60, 240, 60, 240, 
    360, 48, 2400, 480, 180, 24, 480, 240, 240, 480, 48, 2160, 2160, 240, 48, 
    0, 90, 2160, 2160, 240, 240, 120, 120, 72, 240, 72, 24, 240, 240, 60, 
    120, 240, 72, 120, 2160, 24, 2160, 90, 72, 24, 24, 240, 240, 240, 0, 72, 
    0, 2160, 60, 2400, 90, 240, 480, 90, 240, 72, 24, 120, -1, 2160, 480, 0 ;

 VRNXI = 720, 480, 240, 720, 240, 720, 600, 1200, 3600, 240, 720, 240, 720, 
    480, 480, 1200, 3600, 480, 920, 240, 720, 240, 480, 720, 1200, 3000, 
    3000, 480, 1200, 0, 650, 3600, 2880, 480, 480, 600, 720, 720, 480, 720, 
    720, 480, 480, 720, 600, 240, 720, 600, 2880, 24, 2880, 720, 720, 24, 24, 
    480, 480, 240, 0, 720, 0, 2880, 720, 3600, 720, 480, 480, 720, 480, 720, 
    960, 600, -1, 2880, 480, 0 ;

 WDLF = 5, 15, 4, 5, 12.5, 1, 1, 5, 4, 15, 1, 5, 5, 4, 15, 1, 4, 12.5, 4, 
    12.5, 2, 1, 4, 15, 2.5, 4, 4, 4, 2.5, 15, 4, 4, 4, 2, 4, 1, 5, 1, 15, 1, 
    5, 4, 15, 5, 1, 4, 1, 1, 1, 12.5, 4, 4, 2.5, 15, 12.5, 4, 4, 4, 15, 2.5, 
    15, 4, 2.5, 4, 1, 5, 4, 1, 4, 1, 1, 1, 15, 1, 12.5, 15 ;

 PB = 0.1, 0.33, 100, 0.1, 0.1, 1, 10, 0.1, 1, 0.33, 1, 0.33, 0.1, 1, 0.33, 
    1, 1, 0.2, 10, 0.1, 0.2, 1, 1, 0.2, 0.1, 10, 10, 1, 0.1, 0.1, 1, 10, 10, 
    0.33, 1, 10, 0.1, 1, 0.33, 1, 0.1, 1, 0.33, 0.1, 1, 100, 1, 10, 10, 0.1, 
    10, 10, 0.1, 0.1, 0.1, 1, 100, 0.1, 0.1, 0.1, 0.1, 10, 0.1, 1, 1, 0.33, 
    100, 1, 1, 1, 1, 1, 0.1, 10, 0.2, 0.1 ;

 GROUPX = 6.5, 9, 12, 6.5, 17, 6.5, 9, 5, 8, 9, 6.5, 9, 6.5, 9, 9, 5, 21, 8, 
    10, 14, 8, 8, 8, 6, 5, 8, 8, 9, 5, 8.5, 9, 10, 8, 8, 8, 7.5, 8, 7, 9, 9, 
    6.5, 9, 9, 5, 5, 12, 7, 9, 9, 19, 12, 9.5, 7, 9, 19, 8, 11, 9, 8.5, 7, 
    8.5, 11, 6.5, 21, 9, 9, 12, 9, 8, 9, 5, 9, 14, 9, 8, 8.5 ;

 XTLI = 2.5, 2.5, 2.5, 2.5, 5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 
    2.5, 2.5, 2.5, 3, 2.5, 4, 3, 2.5, 2.5, 3, 2.5, 2.5, 2.5, 2.5, 2.5, 3, 
    2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 
    2.5, 2.5, 2.5, 2.5, 2.5, 5, 2.5, 2.5, 2.5, 3, 5, 2.5, 2.5, 2.5, 3, 2.5, 
    3, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 3, 2.5, 3, 3 ;

 XDL = -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 17, 
    -1, -1, -1, -1, -1, -1, -1, -1, 17, 17, -1, -1, -1, -1, -1, 17, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 17, -1, -1, -1, -1, -1, -1, -1, 
    -1, 10, -1, -1, -1 ;

 XPPD = 0.5, 0.5, 2, 0.5, 0.25, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0, 4, 0.5, 0.25, 4, 0.5, 0.5, 4, 0.5, 0, 0, 0.5, 0.5, 0.25, 
    0.5, 1, 0, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 2, 
    0.5, 0.5, 1, 0.25, 1, 0.5, 0.5, 0.25, 0.25, 0.5, 2, 1, 0.25, 0.5, 0.25, 
    1, 0.5, 0, 0.5, 0.5, 2, 0.5, 0.5, 0.5, 0.5, 0.5, 0.15, 1, 4, 0.25 ;

 SLA1 = 0.00333, 0.00333, 0.009, 0.003, 0.015, 0.00167, 0.0125, 0.00333, 
    0.0125, 0.00667, 0.00167, 0.00667, 0.00333, 0.0135, 0.00333, 0.00167, 
    0.009, 0.003, 0.00667, 0.01, 0.003, 0.0333, 0.009, 0.00333, 0.009, 
    0.00667, 0.007, 0.009, 0.00667, 0.00667, 0.009, 0.0083, 0.00667, 0.033, 
    0.009, 0.01, 0.01, 0.00167, 0.00333, 0.00167, 0.00333, 0.0135, 0.00333, 
    0.00333, 0.0033, 0.009, 0.00167, 0.01, 0.01, 0.009, 0.01, 0.00667, 0.009, 
    0.00375, 0.009, 0.009, 0.009, 0.009, 0.00667, 0.009, 0.00667, 0.00667, 
    0.008, 0.009, 0.00333, 0.00333, 0.033, 0.00333, 0.009, 0.00167, 0.00167, 
    0.0033, 0.01, 0.01, 0.003, 0.00667 ;

 SSL1 = 0.125, 0.125, 0.125, 0.125, 0.125, 0.0125, 0.01, 0.125, 0.05, 0.2, 
    0.0125, 0.2, 0.125, 0.125, 0.125, 0.015, 0.015, 0.125, 0.015, 0.125, 
    0.125, 0.01, 0.015, 0.125, 0.0125, 0.015, 0.015, 0.015, 0.0125, 0.2, 
    0.015, 0.05, 0.015, 0.01, 0.125, 0.01, 0.125, 0.015, 0.125, 0.015, 0.125, 
    0.125, 0.125, 0.125, 0.01, 0.125, 0.015, 0.01, 0.01, 0.125, 0.01, 0.015, 
    0.0125, 0.125, 0.125, 0.125, 0.015, 0.015, 0.2, 0.0125, 0.2, 0.015, 
    0.0125, 0.125, 0.015, 0.125, 0.01, 0.015, 0.125, 0.015, 0.0125, 0.01, 
    0.5, 0.01, 0.125, 0.2 ;

 SNL1 = 0.15, 0.15, 0.15, 0.15, 0.25, 0.015, 0.075, 0.15, 0.6, 0.2, 0.015, 
    0.2, 0.15, 0.15, 0.15, 0.015, 0.15, 0.15, 0.15, 0.25, 0.15, 0.075, 0.15, 
    0.15, 0.015, 0.15, 0.15, 0.15, 0.015, 0.2, 0.15, 0.6, 0.15, 0.075, 0.15, 
    0.015, 0.15, 0.015, 0.15, 0.015, 0.15, 0.15, 0.15, 0.15, 0.075, 0.15, 
    0.015, 0.075, 0.075, 0.15, 0.075, 0.15, 0.015, 0.15, 0.15, 0.15, 0.15, 
    0.15, 0.2, 0.015, 0.2, 0.15, 0.015, 0.15, 0.015, 0.15, 0.075, 0.015, 
    0.15, 0.015, 0.015, 0.075, 0.3, 0.075, 0.15, 0.2 ;

 CLASS =
  0, 0, 0.5, 0.5,
  0, 0, 0.5, 0.5,
  0.25, 0.25, 0.25, 0.25,
  0, 0, 0.5, 0.5,
  0, 0, 0.5, 0.5,
  0.25, 0.25, 0.25, 0.25,
  0.25, 0.25, 0.25, 0.25,
  0, 0, 0.5, 0.5,
  0.25, 0.25, 0.25, 0.25,
  0, 0, 0.5, 0.5,
  0.25, 0.25, 0.25, 0.25,
  0.25, 0.25, 0.25, 0.25,
  0, 0, 0.5, 0.5,
  0.25, 0.25, 0.25, 0.25,
  0, 0, 0.5, 0.5,
  0.25, 0.25, 0.25, 0.25,
  0.25, 0.25, 0.25, 0.25,
  0, 0, 0.5, 0.5,
  0.25, 0.25, 0.25, 0.25,
  0.25, 0.25, 0.25, 0.25,
  0.25, 0.25, 0.25, 0.25,
  0.25, 0.25, 0.25, 0.25,
  0.25, 0.25, 0.25, 0.25,
  0, 0, 0.5, 0.5,
  0.25, 0.25, 0.25, 0.25,
  0.25, 0.25, 0.25, 0.25,
  0.25, 0.25, 0.25, 0.25,
  0.25, 0.25, 0.25, 0.25,
  0.25, 0.25, 0.25, 0.25,
  0, 0, 0.5, 0.5,
  0.25, 0.25, 0.25, 0.25,
  0.25, 0.25, 0.25, 0.25,
  0.25, 0.25, 0.25, 0.25,
  0.25, 0.25, 0.25, 0.25,
  0.25, 0.25, 0.25, 0.25,
  0.25, 0.25, 0.25, 0.25,
  0, 0, 0.5, 0.5,
  0.25, 0.25, 0.25, 0.25,
  0, 0, 0.5, 0.5,
  0.25, 0.25, 0.25, 0.25,
  0, 0, 0.5, 0.5,
  0.25, 0.25, 0.25, 0.25,
  0, 0, 0.5, 0.5,
  0, 0, 0.5, 0.5,
  0.25, 0.25, 0.25, 0.25,
  0.25, 0.25, 0.25, 0.25,
  0.25, 0.25, 0.25, 0.25,
  0.25, 0.25, 0.25, 0.25,
  0.25, 0.25, 0.25, 0.25,
  0, 0, 0.5, 0.5,
  0.25, 0.25, 0.25, 0.25,
  0.25, 0.25, 0.25, 0.25,
  0.25, 0.25, 0.25, 0.25,
  0, 0, 0.5, 0.5,
  0.25, 0.25, 0.25, 0.25,
  0.25, 0.25, 0.25, 0.25,
  0.25, 0.25, 0.25, 0.25,
  0.25, 0.25, 0.25, 0.25,
  0, 0, 0.5, 0.5,
  0.25, 0.25, 0.25, 0.25,
  0, 0, 0.5, 0.5,
  0.25, 0.25, 0.25, 0.25,
  0.25, 0.25, 0.25, 0.25,
  0.25, 0.25, 0.25, 0.25,
  0.25, 0.25, 0.25, 0.25,
  0.25, 0.25, 0.25, 0.25,
  0.25, 0.25, 0.25, 0.25,
  0.25, 0.25, 0.25, 0.25,
  0.25, 0.25, 0.25, 0.25,
  0.25, 0.25, 0.25, 0.25,
  0.25, 0.25, 0.25, 0.25,
  0.25, 0.25, 0.25, 0.25,
  0, 0, 0.7, 0.3,
  0.25, 0.25, 0.25, 0.25,
  0, 0, 0.5, 0.5,
  0, 0, 0.5, 0.5 ;

 CFI = 0.9, 1, 1, 0.9, 0.9, 1, 0.5, 0.95, 0.875, 1, 1, 1, 0.9, 1, 1, 1, 0.65, 
    0.8, 0.45, 0.9, 0.9, 0.65, 0.7, 1, 0.65, 0.475, 0.75, 0.65, 0.45, 0.95, 
    0.65, 0.5, 0.45, 0.875, 1, 0.4, 0.9, 1, 1, 1, 0.9, 1, 1, 1, 1, 1, 1, 
    0.45, 0.5, 0.95, 0.5, 0.475, 0.667, 0.95, 0.95, 1, 0.65, 0.7, 0.95, 0.65, 
    0.95, 0.45, 0.475, 1, 1, 1, 0.75, 1, 1, 1, 1, 1, 0.95, 0.7, 0.8, 0.95 ;

 ANGBR = 90, 90, 90, 90, 90, 90, 90, 90, 45, 90, 90, 90, 90, 90, 90, 90, 90, 
    90, 90, 45, 40, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 
    90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 
    90, 45, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 
    90, 60, 90, 90, 90 ;

 ANGSH = 90, 90, 45, 90, 90, 0, 0, 90, 0, 90, 0, 45, 90, 45, 90, 45, 0, 90, 
    0, 45, 45, 45, 0, 90, 0, 0, 0, 45, 0, 90, 0, 0, 0, 0, 45, 0, 90, 45, 90, 
    45, 90, 45, 90, 90, 45, 45, 45, 0, 0, 90, 0, 0, 0, 90, 45, 45, 0, 0, 90, 
    0, 90, 0, 0, 45, 45, 90, 0, 45, 45, 45, 0, 45, 70, 0, 90, 90 ;

 STMX = 5, 3, 1, 5, 5, 10, 0.05, 5, 0.5, 1, 10, 2, 5, 0.5, 3, 10, 1, 7.5, 
    0.1, 4, 7.5, 0.25, 0.5, 7.5, 1, 0.1, 0.1, 0.5, 1, 8, 0.5, 0.1, 0.1, 1, 
    0.5, 0.05, 5, 10, 3, 10, 5, 0.5, 3, 5, 5, 1, 10, 0.05, 0.05, 4, 0.05, 
    0.1, 1, 15, 3, 0.5, 1, 1, 8, 1, 8, 0.1, 1, 1, 10, 3, 0.5, 10, 0.5, 10, 
    10, 5, 120, 0.05, 7.5, 8 ;

 SDMX = 5, 6, 1, 5, 3, 10, 0.1, 5, 1, 6, 10, 6, 5, 1, 6, 10, 1, 6, 0.1, 2, 6, 
    1, 1, 6, 1, 0.1, 50, 1, 1, 6, 1, 0.1, 0.1, 6, 1, 0.1, 5, 10, 6, 10, 5, 1, 
    6, 5, 10, 1, 10, 0.1, 0.1, 3, 0.1, 0.1, 1, 6, 3, 1, 1, 1, 6, 1, 6, 0.1, 
    1, 1, 10, 6, 1, 10, 1, 10, 10, 10, 1, 50, 6, 6 ;

 GRMX = 0.005, 0.01, 0.1, 0.005, 0.2, 0.001, 10, 0.005, 0.1, 0.002, 0.001, 
    0.001, 0.005, 0.1, 0.01, 0.001, 0.1, 0.02, 10, 0.2, 0.02, 0.1, 0.1, 0.02, 
    0.1, 10, 0.02, 0.1, 0.1, 0.02, 0.1, 10, 10, 0.01, 0.1, 10, 0.005, 0.001, 
    0.01, 0.001, 0.005, 0.1, 0.01, 0.005, 0.0001, 0.1, 0.001, 10, 10, 0.2, 
    10, 10, 0.1, 0.02, 0.2, 0.1, 0.1, 0.1, 0.02, 0.1, 0.02, 10, 0.1, 0.1, 
    0.001, 0.01, 0.1, 0.001, 0.1, 0.001, 0.001, 0.0001, 0.01, 0.005, 0.02, 
    0.02 ;

 GRDM = 0.005, 0.01, 1, 0.005, 0.15, 0.001, 10, 0.005, 10, 0.002, 0.001, 
    0.001, 0.005, 1, 0.01, 0.001, 10, 0.02, 10, 0.08, 0.02, 10, 10, 0.02, 1, 
    10, 0.02, 10, 1, 0.02, 10, 10, 10, 0.1, 1, 10, 0.005, 0.001, 0.01, 0.001, 
    0.005, 1, 0.01, 0.5, 0.0001, 1, 0.001, 10, 10, 0.4, 10, 10, 1, 0.04, 0.4, 
    1, 10, 10, 0.02, 1, 0.02, 10, 1, 1, 0.001, 0.01, 10, 0.001, 1, 0.001, 
    0.001, 0.0001, 0.01, 0.005, 0.02, 0.02 ;

 GFILL = 1.25e-05, 2e-05, 0.0002, 1.25e-05, 0.0005, 2.5e-06, 0.02, 1.25e-05, 
    0.0002, 2e-05, 2.5e-06, 2e-05, 1.25e-05, 0.0002, 2e-05, 2.5e-06, 0.0002, 
    5e-05, 0.02, 0.0005, 5e-05, 0.0002, 0.0002, 5e-05, 0.0002, 0.02, 0.02, 
    0.0002, 0.0002, 4e-05, 0.0002, 0.02, 0.02, 2e-05, 0.0002, 0.02, 1.25e-05, 
    2.5e-06, 2e-05, 2.5e-06, 1.25e-05, 0.0002, 2e-05, 1.25e-05, 2.5e-06, 
    0.0002, 2.5e-06, 0.02, 0.02, 0.0005, 0.02, 0.02, 0.0002, 5e-05, 0.0005, 
    0.0002, 0.0002, 0.0002, 4e-05, 0.0002, 4e-05, 0.02, 0.0002, 0.0002, 
    2.5e-06, 2e-05, 0.0002, 2.5e-06, 0.0002, 2.5e-06, 2.5e-06, 2.5e-06, 
    5e-05, 0.02, 5e-05, 4e-05 ;

 WTSTDI = 0, 0, 0, 0, 0, 0, 1000, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4000, 0, 1000, 
    0, 0, 5000, 5000, 0, 100, 5000, 5000, 1000, 100, 0, 5000, 0, 5000, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1000, 5000, 0, 0, 1000, 100, 0, 0, 0, 
    0, 0, 0, 100, 0, 0, 100, 1000, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5000, 0, 0 ;

 RRAD1M = 0.0001, 0.0001, 0.0005, 0.0001, 0.00033, 0.0001, 0.001, 0.0001, 
    0.001, 0.0001, 0.0001, 0.00025, 0.0001, 0.0005, 0.0001, 0.0001, 0.001, 
    0.0002, 0.001, 0.00033, 0.0002, 0.001, 0.001, 0.0002, 0.0005, 0.001, 
    0.001, 0.001, 0.0005, 0.0002, 0.001, 0.001, 0.001, 0.0002, 0.0005, 0.001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0005, 0.0001, 0.0001, 0.0001, 
    0.0005, 0.0001, 0.001, 0.001, 0.0005, 0.001, 0.001, 0.0005, 0.0002, 
    0.00025, 0.0005, 0.001, 0.001, 0.0002, 0.0005, 0.0002, 0.001, 0.00025, 
    0.0005, 0.0001, 0.00025, 0.001, 0.0001, 0.0005, 0.0001, 0.0001, 0.0001, 
    0.0002, 0.0015, 0.0002, 0.0002 ;

 RRAD2M = 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 5e-06, 0.0001, 0.0001, 
    0.0002, 0.0001, 5e-06, 0.0001, 0.0001, 0.0001, 0.0001, 5e-06, 0.0002, 
    0.0001, 0.0002, 6e-06, 0.0001, 0.0001, 0.0002, 0.0001, 0.0001, 0.0002, 
    0.0002, 0.0002, 0.0001, 0.0001, 0.0002, 0.0002, 0.0002, 0.0001, 0.0001, 
    0.0001, 0.0001, 5e-06, 0.0001, 5e-06, 0.0001, 0.0001, 0.0001, 0.0001, 
    5e-06, 0.0001, 5e-06, 0.0001, 0.0001, 0.0001, 0.0001, 0.0002, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0002, 0.0002, 0.0001, 0.0001, 0.0001, 0.0002, 
    0.0001, 0.0001, 5e-06, 0.0001, 0.0001, 5e-06, 0.0001, 5e-06, 5e-06, 
    5e-06, 0.0001, 0.0001, 0.0001, 0.0001 ;

 PORT = 0.05, 0.33, 0.05, 0.45, 0.2, 0, 0.1, 0.05, 0.1, 0.2, 0, 0.2, 0.05, 
    0.25, 0.33, 0, 0.05, 0.2, 0.005, 0.15, 0.2, 0.1, 0.1, 0.2, 0.05, 0.1, 
    0.01, 0.1, 0.05, 0.2, 0.05, 0.25, 0.1, 0.1, 0.2, 0, 0.35, 0, 0.1, 0, 
    0.05, 0.25, 0.1, 0.67, 0, 0.05, 0, 0, 0.1, 0.175, 0.1, 0.1, 0.33, 0.1, 
    0.2, 0.2, 0.05, 0.2, 0.2, 0.05, 0.2, 0.05, 0.05, 0.05, 0.01, 0.2, 0.1, 
    0.01, 0.2, 0, 0, 0, 0.4, 0.1, 0.2, 0.2 ;

 PR = 0.1, 0.1, 0.2, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 
    0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 
    0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 
    0.1, 0.1, 0.1, 0.2, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 
    0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.05, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 
    0.1, 0.1, 0.1, 0.1, 0.1, 0.1 ;

 RSRR = 10000, 10000, 10000, 500000, 10000, 10000, 10000, 10000, 10000, 
    10000, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 500000, 
    40000, 20000, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 
    10000, 10000, 10000, 10000, 10000, 10000, 10000, 500000, 10000, 10000, 
    10000, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 
    10000, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 
    10000, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 10000, 
    10000, 10000, 10000, 2500, 10000, 10000, 10000 ;

 RSRA = 4e+09, 4e+09, 4e+09, 1000000, 5e+07, 4e+09, 1e+10, 4e+09, 4e+09, 
    1e+09, 4e+09, 1e+09, 4e+09, 4e+09, 4e+09, 4e+09, 4e+09, 2e+08, 1000, 
    1e+08, 2e+08, 1e+09, 4e+09, 4e+08, 4e+09, 4e+10, 2e+09, 4e+09, 4e+10, 
    1e+09, 4e+09, 4e+09, 4e+10, 1e+09, 4e+09, 1e+10, 1000000, 4e+09, 4e+09, 
    4e+09, 4e+09, 4e+09, 4e+09, 4e+09, 1e+10, 4e+09, 4e+09, 1e+10, 1e+10, 
    4e+08, 1e+10, 4e+10, 4e+09, 4e+08, 4e+08, 4e+09, 4e+09, 4e+09, 1e+09, 
    4e+09, 1e+09, 4e+10, 4e+10, 4e+09, 4e+09, 4e+09, 1e+09, 4e+09, 4e+09, 
    4e+09, 4e+09, 1e+10, 4e+08, 1e+10, 2e+08, 1e+09 ;

 PTSHT = 0.05, 0.05, 0.01, 0.04, 0.03, 0.001, 0.01, 0.01, 0.0075, 0.05, 
    0.001, 0.025, 0.05, 0.01, 0.05, 0.0001, 0.01, 0.05, 0.01, 0.008, 0.05, 
    0.01, 0.01, 0.05, 0.01, 0.01, 0.1, 0.01, 0.01, 0.025, 0.01, 0.00375, 
    0.01, 0.025, 0.01, 0.01, 0.05, 0.01, 0.05, 0.01, 0.05, 0.01, 0.05, 0.05, 
    0.01, 0.01, 0.0001, 0.01, 0.01, 0.05, 0.01, 0.01, 0.01, 0.05, 0.05, 0.01, 
    0.01, 0.01, 0.025, 0.01, 0.025, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.05, 0.01, 0.025, 0.01, 0.05, 0.025 ;

 RTFQ = 250, 250, 250, 1200, 500, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 40, 400, 250, 250, 250, 250, 250, 250, 300, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 300, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 
    250, 250, 800, 500, 250, 250 ;

 UPMXZH = 0.005, 0.005, 0.005, 0.005, 0.025, 0, 0.0025, 0.005, 0.005, 0.01, 
    0, 0.01, 0.005, 0.005, 0.005, 5e-05, 0.005, 0.025, 0.005, 0.03, 0.025, 
    0.0025, 0.005, 0.025, 0.005, 0.005, 0.005, 0.005, 0.005, 0.01, 0.005, 
    0.005, 0.005, 0.0025, 0.005, 0.0025, 0.005, 5e-05, 0.005, 5e-05, 0.005, 
    0.005, 0.005, 0.005, 5e-05, 0.005, 5e-05, 0.0025, 0.0025, 0.025, 0.0025, 
    0.005, 0.005, 0.025, 0.025, 0.005, 0.005, 0.0005, 0.01, 0.005, 0.01, 
    0.005, 0.005, 0.005, 0.0005, 0.005, 0.0025, 0.0005, 0.005, 5e-05, 0.005, 
    3.3e-05, 0.025, 0.0025, 0.025, 0.01 ;

 UPKMZH = 0.4, 0.4, 0.4, 0.4, 5, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 
    0.4, 0.4, 0.4, 4, 0.4, 4, 4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 
    0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 
    0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 
    0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 
    0.4, 0.4, 4, 0.4 ;

 UPMNZH = 0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 
    0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 
    0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 
    0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 
    0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 
    0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 
    0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 
    0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 
    0.0125, 0.0125, 0.0125, 0.0125, 0.0125 ;

 UPMXZO = 0.005, 0.005, 0.005, 0.005, 0.1, 0, 0.0025, 0.005, 0.005, 0.01, 0, 
    0.01, 0.005, 0.005, 0.005, 5e-05, 0.005, 0.025, 0.005, 0.1, 0.025, 
    0.0025, 0.005, 0.025, 0.005, 0.005, 0.005, 0.005, 0.005, 0.01, 0.005, 
    0.005, 0.005, 0.0025, 0.005, 0.0025, 0.005, 5e-05, 0.005, 5e-05, 0.005, 
    0.005, 0.005, 0.005, 5e-05, 0.005, 5e-05, 0.0025, 0.0025, 0.025, 0.0025, 
    0.005, 0.005, 0.025, 0.025, 0.005, 0.005, 0.0005, 0.01, 0.005, 0.01, 
    0.005, 0.005, 0.005, 0.0005, 0.005, 0.0025, 0.0005, 0.005, 5e-05, 0.005, 
    3.3e-05, 0.025, 0.0025, 0.025, 0.01 ;

 UPKMZO = 0.35, 0.35, 0.35, 0.35, 10, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 
    0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 6, 0.35, 15, 6, 0.35, 0.35, 0.35, 
    0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 
    0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 
    0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 
    0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 
    0.35, 0.35, 6, 0.35 ;

 UPMNZO = 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 
    0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 
    0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 
    0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 
    0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 
    0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 
    0.03, 0.03, 0.03, 0.03, 0.03 ;

 UPMXPO = 0.001, 0.001, 0.001, 0.001, 0.005, 0.001, 0.0025, 0.001, 0.001, 
    0.01, 0.001, 0.01, 0.001, 0.001, 0.001, 0.001, 0.0005, 0.005, 0.001, 
    0.005, 0.005, 0.0025, 0.001, 0.005, 0.001, 0.001, 0.001, 0.001, 0.001, 
    0.01, 0.001, 0.001, 0.001, 0.0025, 0.001, 0.0025, 0.001, 0.001, 0.001, 
    0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.0025, 0.0025, 
    0.005, 0.0025, 0.001, 0.001, 0.005, 0.005, 0.001, 0.001, 0.001, 0.01, 
    0.001, 0.01, 0.001, 0.001, 0.0005, 0.001, 0.001, 0.0025, 0.001, 0.001, 
    0.001, 0.001, 0.001, 0.025, 0.0025, 0.005, 0.01 ;

 UPKMPO = 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 
    0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 
    0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 
    0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 
    0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 
    0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 
    0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 
    0.075, 0.075, 0.075, 0.075, 0.075, 0.075, 0.075 ;

 UPMNPO = 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002 ;

 OSMO = -1.25, -1.25, -1.25, -1.25, -1.25, -1.25, -1.5, -1.25, -1.25, -1.25, 
    -1.25, -1.25, -1.25, -1.25, -1.25, -1.25, -1.5, -1.25, -1.25, -1.5, 
    -1.25, -1.25, -1.25, -1.25, -1.25, -1.25, -1.25, -1.25, -1.25, -1.25, 
    -1.25, -1.25, -1.25, -1.25, -1.25, -1.25, -1.25, -1.25, -1.25, -1.25, 
    -1.25, -1.25, -1.25, -1.25, -1.25, -1.25, -1.25, -1.25, -1.25, -1.25, 
    -1.5, -1.25, -1.25, -1.25, -1.25, -1.25, -1.25, -1.25, -1.25, -1.25, 
    -1.25, -1.25, -1.25, -1.5, -1.25, -1.25, -1.25, -1.25, -1.25, -2.5, 
    -1.25, -1.25, -2, -1.25, -1.25, -1.25 ;

 RCS = 0.2, 0.2, 0.2, 0.125, 0.2, 100, 0.2, 0.2, 0.2, 0.2, 100, 0.2, 0.2, 
    0.2, 0.2, 100, 0.2, 0.2, 0.2, 0.2, 0.2, 0.2, 0.2, 0.2, 0.2, 0.2, 0.2, 
    0.2, 0.2, 0.2, 0.2, 0.2, 0.2, 0.2, 0.2, 0.2, 0.2, 100, 0.2, 0, 0.2, 0.2, 
    0.2, 0.2, 100, 0.2, 100, 0.2, 0.2, 0.2, 0.2, 0.2, 0.2, 0.2, 0.2, 0.2, 
    0.2, 0.2, 0.2, 0.2, 0.2, 0.2, 0.2, 0.2, 0, 0.2, 0.2, 100, 0.2, 100, 100, 
    100, 0.125, 0.2, 0.2, 0.2 ;

 RSMX = 2500, 5000, 2500, 2500, 5000, 500, 5000, 2500, 5000, 5000, 500, 5000, 
    2500, 2500, 5000, 500, 5000, 2500, 2500, 5000, 2500, 2500, 2500, 2500, 
    2500, 2500, 3500, 2000, 2500, 2000, 2000, 5000, 2500, 5000, 2500, 2500, 
    2500, 150, 5000, 150, 2500, 2500, 5000, 2500, 200, 2500, 500, 2500, 5000, 
    5000, 5000, 2500, 2500, 2000, 5000, 2500, 5000, 2500, 2000, 2500, 2000, 
    2500, 2500, 5000, 150, 5000, 5000, 150, 2500, 600, 150, 600, 2000, 2000, 
    2500, 2000 ;

 DMLF = 0.72, 0.72, 0.72, 0.72, 0.72, 0.76, 0.76, 0.72, 0.72, 0.72, 0.76, 
    0.72, 0.72, 0.72, 0.72, 0.76, 0.72, 0.72, 0.76, 0.67, 0.72, 0.72, 0.72, 
    0.72, 0.72, 0.76, 0.76, 0.72, 0.76, 0.72, 0.72, 0.76, 0.76, 0.72, 0.72, 
    0.76, 0.72, 0.76, 0.72, 0.76, 0.72, 0.72, 0.72, 0.72, 0.76, 0.72, 0.76, 
    0.76, 0.76, 0.72, 0.76, 0.76, 0.72, 0.72, 0.72, 0.72, 0.72, 0.72, 0.72, 
    0.72, 0.72, 0.76, 0.76, 0.72, 0.76, 0.72, 0.72, 0.76, 0.72, 0.76, 0.76, 
    0.76, 0.72, 0.76, 0.72, 0.72 ;

 DMSHE = 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 
    0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 
    0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 
    0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 
    0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 
    0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 
    0.76, 0.76, 0.76, 0.76, 0.76 ;

 DMSTK = 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 
    0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 
    0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 
    0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 
    0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 
    0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8 ;

 DMRSV = 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 
    0.67, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.67, 0.88, 0.88, 0.88, 
    0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 
    0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 
    0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.67, 0.88, 0.88, 0.88, 0.88, 
    0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.67, 0.88, 0.88, 0.88, 0.88, 0.88, 
    0.88, 0.88, 0.88, 0.88, 0.88 ;

 DMHSK = 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 
    0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 
    0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 
    0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 
    0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 
    0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 
    0.76, 0.76, 0.76, 0.76, 0.76 ;

 DMEAR = 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 
    0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 
    0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 
    0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 
    0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 
    0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 
    0.76, 0.76, 0.76, 0.76, 0.76 ;

 DMGR = 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 
    0.67, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.67, 0.88, 0.88, 0.88, 
    0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 
    0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 
    0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.67, 0.88, 0.88, 0.88, 0.88, 
    0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.67, 0.88, 0.88, 0.88, 0.88, 0.88, 
    0.88, 0.88, 0.88, 0.88, 0.88 ;

 DMRT = 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 
    0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 
    0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 
    0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 
    0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 
    0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 
    0.76, 0.76, 0.76, 0.76, 0.76 ;

 DMND = 0.72, 0.72, 0.72, 0.72, 0.72, 0.72, 0.5, 0.72, 0.72, 0.5, 0.72, 0.5, 
    0.72, 0.72, 0.72, 0.72, 0.72, 0.72, 0.72, 0.67, 0.72, 0.5, 0.72, 0.72, 
    0.72, 0.72, 0.72, 0.72, 0.72, 0.5, 0.72, 0.72, 0.72, 0.5, 0.72, 0.5, 
    0.72, 0.72, 0.72, 0.72, 0.72, 0.72, 0.72, 0.72, 0.5, 0.72, 0.72, 0.5, 
    0.5, 0.72, 0.5, 0.72, 0.72, 0.72, 0.67, 0.72, 0.72, 0.72, 0.5, 0.72, 0.5, 
    0.72, 0.72, 0.72, 0.72, 0.67, 0.5, 0.72, 0.72, 0.72, 0.72, 0.5, 0.6, 0.5, 
    0.72, 0.5 ;

 CNWR = 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 
    2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 
    2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 
    2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 
    2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 
    2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 2.15, 
    2.15, 2.15, 2.15, 2.15, 2.15 ;

 CNWL = 2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 
    2.6, 2.6, 2.6, 3.5, 2.6, 2.6, 3.5, 2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 
    2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 
    2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 
    2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 2.6, 
    2.6, 2.6, 2.6, 2.6, 3.5, 2.6 ;

 CNLF = 0.1, 0.1, 0.1, 0.03, 0.1, 0.04, 0.0333, 0.1, 0.1, 0.1, 0.04, 0.1, 
    0.1, 0.1, 0.1, 0.0333, 0.1, 0.1, 0.0333, 0.15, 0.1, 0.0833, 0.1, 0.1, 
    0.1, 0.04, 0.04, 0.1, 0.0333, 0.1, 0.1, 0.045, 0.0333, 0.0833, 0.1, 
    0.0333, 0.1, 0.0333, 0.1, 0.0333, 0.1, 0.1, 0.1, 0.1, 0.0833, 0.1, 
    0.0333, 0.0333, 0.0333, 0.1, 0.0333, 0.04, 0.1, 0.1, 0.125, 0.1, 0.1, 
    0.1, 0.1, 0.1, 0.1, 0.0333, 0.04, 0.1, 0.04, 0.1, 0.0833, 0.04, 0.1, 
    0.0333, 0.0333, 0.0833, 0.1, 0.0333, 0.1, 0.1 ;

 CNSHE = 0.02, 0.02, 0.02, 0.006, 0.025, 0.02, 0.02, 0.02, 0.025, 0.025, 
    0.02, 0.025, 0.02, 0.02, 0.02, 0.02, 0.02, 0.025, 0.02, 0.0375, 0.025, 
    0.02, 0.02, 0.025, 0.02, 0.02, 0.02, 0.02, 0.02, 0.025, 0.02, 0.02, 0.02, 
    0.025, 0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 
    0.02, 0.02, 0.02, 0.02, 0.025, 0.02, 0.02, 0.02, 0.025, 0.025, 0.02, 
    0.02, 0.025, 0.025, 0.02, 0.025, 0.02, 0.02, 0.02, 0.02, 0.025, 0.02, 
    0.02, 0.02, 0.02, 0.02, 0.02, 0.025, 0.02, 0.025, 0.025 ;

 CNSTK = 0.01, 0.01, 0.004, 0.003, 0.01, 0.01, 0.004, 0.01, 0.004, 0.01, 
    0.01, 0.02, 0.01, 0.004, 0.01, 0.01, 0.004, 0.01, 0.004, 0.02, 0.02, 
    0.004, 0.004, 0.01, 0.004, 0.004, 0.004, 0.004, 0.004, 0.01, 0.004, 
    0.004, 0.004, 0.01, 0.004, 0.004, 0.01, 0.01, 0.01, 0.01, 0.01, 0.004, 
    0.01, 0.01, 0.01, 0.004, 0.01, 0.004, 0.004, 0.01, 0.004, 0.004, 0.004, 
    0.01, 0.02, 0.004, 0.004, 0.004, 0.01, 0.004, 0.01, 0.004, 0.004, 0.004, 
    0.01, 0.02, 0.004, 0.01, 0.004, 0.01, 0.01, 0.01, 0.01, 0.004, 0.01, 0.01 ;

 CNRSV = 0.02, 0.025, 0.04, 0.006, 0.03, 0.02, 0.02, 0.02, 0.02, 0.04, 0.02, 
    0.125, 0.02, 0.02, 0.025, 0.02, 0.02, 0.04, 0.03, 0.125, 0.1, 0.02, 0.02, 
    0.04, 0.02, 0.02, 0.02, 0.02, 0.02, 0.04, 0.04, 0.02, 0.02, 0.04, 0.02, 
    0.02, 0.02, 0.02, 0.025, 0.02, 0.02, 0.02, 0.025, 0.02, 0.02, 0.04, 0.02, 
    0.02, 0.02, 0.03, 0.02, 0.03, 0.02, 0.04, 0.1, 0.02, 0.04, 0.02, 0.04, 
    0.02, 0.04, 0.02, 0.02, 0.04, 0.02, 0.125, 0.04, 0.02, 0.02, 0.02, 0.02, 
    0.02, 0.04, 0.02, 0.04, 0.04 ;

 CNHSK = 0.02, 0.02, 0.02, 0.006, 0.02, 0.02, 0.02, 0.02, 0.02, 0.025, 0.02, 
    0.025, 0.02, 0.02, 0.02, 0.02, 0.02, 0.025, 0.02, 0.025, 0.025, 0.02, 
    0.02, 0.025, 0.02, 0.02, 0.02, 0.02, 0.02, 0.025, 0.02, 0.02, 0.02, 
    0.025, 0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 
    0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 0.025, 0.025, 0.02, 0.02, 
    0.02, 0.025, 0.02, 0.025, 0.02, 0.02, 0.02, 0.02, 0.025, 0.02, 0.02, 
    0.02, 0.02, 0.02, 0.02, 0.025, 0.02, 0.025, 0.025 ;

 CNEAR = 0.02, 0.02, 0.02, 0.006, 0.02, 0.02, 0.02, 0.02, 0.02, 0.025, 0.02, 
    0.025, 0.02, 0.02, 0.02, 0.02, 0.02, 0.025, 0.02, 0.025, 0.025, 0.02, 
    0.02, 0.025, 0.02, 0.02, 0.02, 0.02, 0.02, 0.025, 0.02, 0.02, 0.02, 
    0.025, 0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 
    0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 0.025, 0.025, 0.02, 0.02, 
    0.02, 0.025, 0.02, 0.025, 0.02, 0.02, 0.02, 0.02, 0.025, 0.02, 0.02, 
    0.02, 0.02, 0.02, 0.02, 0.025, 0.02, 0.025, 0.025 ;

 CNGR = 0.04, 0.033, 0.04, 0.012, 0.0375, 0.04, 0.04, 0.04, 0.02, 0.055, 
    0.04, 0.15, 0.04, 0.04, 0.033, 0.04, 0.04, 0.055, 0.04, 0.15, 0.125, 
    0.04, 0.04, 0.055, 0.04, 0.04, 0.04, 0.04, 0.04, 0.055, 0.04, 0.02, 0.04, 
    0.055, 0.04, 0.04, 0.04, 0.04, 0.033, 0.04, 0.04, 0.04, 0.033, 0.04, 
    0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.02, 0.04, 0.04, 0.055, 0.14, 0.04, 
    0.04, 0.02, 0.055, 0.04, 0.055, 0.02, 0.04, 0.05, 0.04, 0.15, 0.04, 0.04, 
    0.04, 0.04, 0.04, 0.04, 0.055, 0.04, 0.055, 0.055 ;

 CNRT = 0.025, 0.025, 0.025, 0.0075, 0.02, 0.02, 0.02, 0.02, 0.02, 0.025, 
    0.02, 0.025, 0.025, 0.02, 0.025, 0.02, 0.02, 0.025, 0.02, 0.025, 0.025, 
    0.02, 0.02, 0.025, 0.02, 0.02, 0.02, 0.02, 0.02, 0.025, 0.02, 0.02, 0.02, 
    0.025, 0.02, 0.02, 0.025, 0.02, 0.025, 0.02, 0.025, 0.02, 0.025, 0.02, 
    0.02, 0.025, 0.02, 0.02, 0.025, 0.025, 0.02, 0.02, 0.02, 0.025, 0.025, 
    0.02, 0.02, 0.025, 0.025, 0.02, 0.025, 0.02, 0.02, 0.02, 0.02, 0.025, 
    0.02, 0.02, 0.02, 0.02, 0.02, 0.02, 0.025, 0.025, 0.025, 0.025 ;

 CNND = 0.1, 0.1, 0.1, 0.03, 0.1, 0.125, 0.125, 0.1, 0.1, 0.1, 0.125, 0.125, 
    0.1, 0.125, 0.1, 0.125, 0.1, 0.1, 0.1, 0.125, 0.125, 0.125, 0.1, 0.1, 
    0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.125, 0.125, 0.125, 0.1, 
    0.125, 0.1, 0.125, 0.1, 0.125, 0.1, 0.1, 0.125, 0.125, 0.125, 0.125, 
    0.125, 0.1, 0.0833, 0.1, 0.1, 0.1, 0.125, 0.125, 0.1, 0.125, 0.1, 0.1, 
    0.1, 0.1, 0.1, 0.1, 0.125, 0.125, 0.1, 0.125, 0.125, 0.125, 0.1, 0.125, 
    0.1, 0.125, 0.1, 0.1 ;

 CPWR = 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 
    40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 
    40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 
    40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 
    40, 40, 40, 40, 40 ;

 CPWL = 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 
    28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 
    28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 
    28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 
    28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 
    28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 28.4, 
    28.4, 28.4, 28.4, 28.4, 28.4 ;

 CPLF = 0.01, 0.01, 0.01, 0.003, 0.01, 0.004, 0.00333, 0.01, 0.01, 0.01, 
    0.004, 0.01, 0.01, 0.01, 0.01, 0.00333, 0.01, 0.01, 0.00333, 0.015, 0.01, 
    0.00833, 0.01, 0.01, 0.01, 0.004, 0.004, 0.01, 0.00333, 0.01, 0.01, 
    0.0045, 0.00333, 0.00833, 0.01, 0.00333, 0.01, 0.00333, 0.01, 0.00333, 
    0.01, 0.01, 0.01, 0.01, 0.00833, 0.01, 0.00333, 0.00333, 0.00333, 0.01, 
    0.00333, 0.004, 0.01, 0.01, 0.0125, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.00333, 0.004, 0.01, 0.004, 0.01, 0.00833, 0.004, 0.01, 0.00333, 
    0.00333, 0.00833, 0.01, 0.00333, 0.01, 0.01 ;

 CPSHE = 0.002, 0.002, 0.002, 0.0006, 0.0025, 0.002, 0.002, 0.002, 0.0025, 
    0.0025, 0.002, 0.0025, 0.002, 0.002, 0.002, 0.002, 0.002, 0.0025, 0.002, 
    0.00375, 0.0025, 0.002, 0.002, 0.0025, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.0025, 0.002, 0.002, 0.002, 0.0025, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.0025, 0.002, 0.002, 0.002, 0.0025, 0.0025, 0.002, 0.002, 0.0025, 
    0.0025, 0.002, 0.0025, 0.002, 0.002, 0.002, 0.002, 0.0025, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.0025, 0.002, 0.0025, 0.0025 ;

 CPSTK = 0.001, 0.001, 0.0004, 0.0003, 0.001, 0.001, 0.0004, 0.001, 0.0004, 
    0.001, 0.001, 0.002, 0.001, 0.0004, 0.001, 0.001, 0.0004, 0.001, 0.0004, 
    0.002, 0.002, 0.0004, 0.0004, 0.001, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.001, 0.0004, 0.0004, 0.0004, 0.001, 0.0004, 0.0004, 0.001, 
    0.001, 0.001, 0.001, 0.001, 0.0004, 0.001, 0.001, 0.001, 0.0004, 0.001, 
    0.0004, 0.0004, 0.001, 0.0004, 0.0004, 0.0004, 0.001, 0.002, 0.0004, 
    0.0004, 0.0004, 0.001, 0.0004, 0.001, 0.0004, 0.0004, 0.0004, 0.001, 
    0.002, 0.0004, 0.001, 0.0004, 0.001, 0.001, 0.001, 0.001, 0.0004, 0.001, 
    0.001 ;

 CPRSV = 0.002, 0.0025, 0.004, 0.0006, 0.003, 0.002, 0.002, 0.002, 0.002, 
    0.004, 0.002, 0.0125, 0.002, 0.002, 0.0025, 0.002, 0.002, 0.004, 0.003, 
    0.0125, 0.01, 0.002, 0.002, 0.004, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.004, 0.004, 0.002, 0.002, 0.004, 0.002, 0.002, 0.002, 0.002, 0.0025, 
    0.002, 0.002, 0.002, 0.0025, 0.002, 0.002, 0.004, 0.002, 0.002, 0.002, 
    0.003, 0.002, 0.003, 0.002, 0.004, 0.01, 0.002, 0.004, 0.002, 0.004, 
    0.002, 0.004, 0.002, 0.002, 0.004, 0.002, 0.0125, 0.004, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.004, 0.002, 0.004, 0.004 ;

 CPHSK = 0.002, 0.002, 0.002, 0.0006, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.0025, 0.002, 0.0025, 0.002, 0.002, 0.002, 0.002, 0.002, 0.0025, 0.002, 
    0.0025, 0.0025, 0.002, 0.002, 0.0025, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.0025, 0.002, 0.002, 0.002, 0.0025, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.0025, 0.0025, 0.002, 0.002, 0.002, 0.0025, 
    0.002, 0.0025, 0.002, 0.002, 0.002, 0.002, 0.0025, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.0025, 0.002, 0.0025, 0.0025 ;

 CPEAR = 0.002, 0.002, 0.002, 0.0006, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.0025, 0.002, 0.0025, 0.002, 0.002, 0.002, 0.002, 0.002, 0.0025, 0.002, 
    0.0025, 0.0025, 0.002, 0.002, 0.0025, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.0025, 0.002, 0.002, 0.002, 0.0025, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.0025, 0.0025, 0.002, 0.002, 0.002, 0.0025, 
    0.002, 0.0025, 0.002, 0.002, 0.002, 0.002, 0.0025, 0.002, 0.002, 0.002, 
    0.002, 0.002, 0.002, 0.0025, 0.002, 0.0025, 0.0025 ;

 CPGR = 0.004, 0.0033, 0.004, 0.0012, 0.00375, 0.004, 0.004, 0.004, 0.002, 
    0.0055, 0.004, 0.015, 0.004, 0.004, 0.0033, 0.004, 0.004, 0.0055, 0.004, 
    0.015, 0.0125, 0.004, 0.004, 0.0055, 0.004, 0.004, 0.004, 0.004, 0.004, 
    0.0055, 0.004, 0.002, 0.004, 0.0055, 0.004, 0.004, 0.004, 0.004, 0.0033, 
    0.004, 0.004, 0.004, 0.0033, 0.004, 0.004, 0.004, 0.004, 0.004, 0.004, 
    0.004, 0.002, 0.004, 0.004, 0.0055, 0.014, 0.004, 0.004, 0.002, 0.0055, 
    0.004, 0.0055, 0.002, 0.004, 0.005, 0.004, 0.015, 0.004, 0.004, 0.004, 
    0.004, 0.004, 0.004, 0.0055, 0.004, 0.0055, 0.0055 ;

 CPRT = 0.0025, 0.0025, 0.0025, 0.00075, 0.002, 0.002, 0.002, 0.002, 0.002, 
    0.0025, 0.002, 0.0025, 0.0025, 0.002, 0.0025, 0.002, 0.002, 0.0025, 
    0.002, 0.0025, 0.0025, 0.002, 0.002, 0.0025, 0.002, 0.002, 0.002, 0.002, 
    0.002, 0.0025, 0.002, 0.002, 0.002, 0.0025, 0.002, 0.002, 0.0025, 0.002, 
    0.0025, 0.002, 0.0025, 0.002, 0.0025, 0.002, 0.002, 0.0025, 0.002, 0.002, 
    0.0025, 0.0025, 0.002, 0.002, 0.002, 0.0025, 0.0025, 0.002, 0.002, 
    0.0025, 0.0025, 0.002, 0.0025, 0.002, 0.002, 0.002, 0.002, 0.0025, 0.002, 
    0.002, 0.002, 0.002, 0.002, 0.002, 0.0025, 0.0025, 0.0025, 0.0025 ;

 CPND = 0.01, 0.01, 0.01, 0.003, 0.01, 0.0125, 0.0125, 0.01, 0.01, 0.01, 
    0.0125, 0.0125, 0.01, 0.0125, 0.01, 0.0125, 0.01, 0.01, 0.01, 0.0125, 
    0.0125, 0.0125, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.0125, 0.0125, 0.0125, 0.01, 0.0125, 0.01, 0.0125, 0.01, 
    0.0125, 0.01, 0.01, 0.0125, 0.0125, 0.0125, 0.0125, 0.0125, 0.01, 
    0.00833, 0.01, 0.01, 0.01, 0.0125, 0.0125, 0.01, 0.0125, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.0125, 0.0125, 0.01, 0.0125, 0.0125, 0.0125, 
    0.01, 0.0125, 0.01, 0.0125, 0.01, 0.01 ;

 ROOTMAGE = 60, 360, 240, 40, 240, 60, 120, 48, 1500, 240, 60, 240, 60, 240, 
    360, 48, 2400, 480, 180, 24, 480, 240, 240, 480, 48, 2160, 2160, 240, 48, 
    0, 90, 2160, 2160, 240, 240, 120, 120, 72, 240, 72, 24, 240, 240, 60, 
    120, 240, 72, 120, 2160, 24, 2160, 90, 72, 24, 24, 240, 240, 240, 0, 72, 
    0, 2160, 60, 2400, 90, 240, 480, 90, 240, 72, 24, 120, -1, 2160, 480, 0 ;

 pfts =
  "gr3s32",
  "gr3s35",
  "bush31",
  "sedg62",
  "maiz31",
  "lich33",
  "jpin43",
  "gr3s61",
  "shru35",
  "brom43",
  "lich32",
  "alfa43",
  "gr3s33",
  "busn32",
  "clvs35",
  "lich61",
  "bdlf11",
  "gr3a35",
  "ndlf43",
  "soyb31",
  "clva35",
  "tasp43",
  "bdlf43",
  "gr3a34",
  "bdlf61",
  "ndlf33",
  "ndlf34",
  "bdlf32",
  "ndlf61",
  "oats43",
  "bdlf33",
  "ndlf35",
  "ndlf32",
  "busn26",
  "busn43",
  "bspr62",
  "gr3s43",
  "moss62",
  "gr3s26",
  "moss43",
  "gr3s62",
  "bush32",
  "gr4s26",
  "sedg61",
  "smos61",
  "busn31",
  "lich62",
  "bspr43",
  "dfir32",
  "maiz33",
  "lpin31",
  "ndld43",
  "bdlw62",
  "swhe33",
  "soyb33",
  "bdln43",
  "bdlf31",
  "bdln32",
  "barl43",
  "bdlf62",
  "swhe43",
  "ndlf31",
  "ndlf62",
  "bush11",
  "moss33",
  "bush26",
  "woak31",
  "moss32",
  "bush43",
  "mosf43",
  "moss61",
  "fmos43",
  "rice34",
  "dfir34",
  "dgra35",
  "woat35" ;

 pfts_short =
  "alfa",
  "barl",
  "bdlf",
  "bdln",
  "bdlw",
  "brom",
  "bspr",
  "fmos",
  "ndlf",
  "ndld",
  "gr3s",
  "gr4s",
  "gr3a",
  "clva",
  "clvs",
  "bush",
  "dfir",
  "busn",
  "lpin",
  "maiz",
  "oats",
  "rice",
  "shru",
  "soyb",
  "swhe",
  "lich",
  "jpin",
  "moss",
  "mosf",
  "smos",
  "sedg",
  "tasp",
  "woak",
  "dgra",
  "woat" ;

 pfts_long =
  "alfalfa crop                            ",
  "barley crop                             ",
  "broadleaf tree (deciduous or evergreen) ",
  "broadleaf tree with N2 fixation         ",
  "broadleaf tree adapted to wetland       ",
  "brome grass                             ",
  "black spruce tree (needle leaf)         ",
  "feather moss (with jack pine)           ",
  "needleleaf tree (evergreen)             ",
  "needleleaf tree (deciduous)             ",
  "C3 grass perennial                      ",
  "C4 grass perennial                      ",
  "C3 grass annual                         ",
  "clover annual crop                      ",
  "clover perennial crop                   ",
  "bush tree                               ",
  "douglas fir tree                        ",
  "bush tree with N2 fixation              ",
  "loblolly pine tree                      ",
  "maize crop                              ",
  "oats crop                               ",
  "rice crop                               ",
  "shrub tree                              ",
  "soybean crop                            ",
  "spring wheat crop                       ",
  "lichen                                  ",
  "jackpine tree                           ",
  "moss (sphagnum)                         ",
  "moss (feathermoss)                      ",
  "moss (sphagnum near sedge)              ",
  "sedge grass                             ",
  "aspen tree                              ",
  "oak tree (upland)                       ",
  "deer grass                              ",
  "wild oats                               " ;

 koppen_clim_no =
  "11",
  "12",
  "13",
  "14",
  "21",
  "22",
  "26",
  "27",
  "31",
  "32",
  "33",
  "34",
  "35",
  "36",
  "37",
  "38",
  "39",
  "41",
  "42",
  "43",
  "44",
  "45",
  "46",
  "47",
  "48",
  "49",
  "50",
  "51",
  "52",
  "61",
  "62" ;

 koppen_clim_short =
  "Af ",
  "Am ",
  "As ",
  "Aw ",
  "BWk",
  "BWh",
  "BSk",
  "BSh",
  "Cfa",
  "Cfb",
  "Cfc",
  "Csa",
  "Csb",
  "Csc",
  "Cwa",
  "Cwb",
  "Cwc",
  "Dfa",
  "Dfb",
  "Dfc",
  "Dfd",
  "Dsa",
  "Dsb",
  "Dsc",
  "Dsd",
  "Dwa",
  "Dwb",
  "Dwc",
  "Dwd",
  "ET ",
  "EF " ;

 koppen_clim_long =
  "Tropical rainforest climate                                     ",
  "Tropical monsoon climate                                        ",
  "Tropical summer-dry climate                                     ",
  "Tropical winter-dry climate                                     ",
  "Cold desert climate                                             ",
  "Hot desert climate                                              ",
  "Cold semi-arid climate                                          ",
  "Hot semi-arid climate                                           ",
  "Humid subtropical climate                                       ",
  "Temperate oceanic climate                                       ",
  "Subpolar oceanic climate                                        ",
  "Hot-summer Mediterranean climate                                ",
  "Warm-summer Mediterranean climate                               ",
  "Cold-summer Mediterranean climate                               ",
  "Monsoon-influenced humid subtropical climate                    ",
  "Subtropical highland climate                                    ",
  "Cold subtropical highland climate                               ",
  "Hot-summer humid continental climate                            ",
  "Warm-summer humid continental climate                           ",
  "Subarctic climate                                               ",
  "Extremely cold subarctic climate                                ",
  "Mediterranean-influenced hot-summer humid continental climate   ",
  "Mediterranean-influenced warm-summer humid continental climate  ",
  "Mediterranean-influenced subarctic climate                      ",
  "Mediterranean-influenced extremely cold subarctic climate       ",
  "Monsoon-influenced hot-summer humid continental climate         ",
  "Monsoon-influenced warm-summer humid continental climate        ",
  "Monsoon-influenced subarctic climate                            ",
  "Monsoon-influenced extremely cold subarctic climate             ",
  "Tundra climate                                                  ",
  "Ice cap climate                                                 " ;
}
