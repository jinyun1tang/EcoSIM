netcdf fatm_hist_GHGs_1750-2023 {
dimensions:
	time = UNLIMITED ; // (3276 currently)
variables:
	float CH4(time) ;
		CH4:long_name = "Atmospheric CH4 concentrations" ;
		CH4:units = "ppbv" ;
	float CO2(time) ;
		CO2:long_name = "Atmospheric CO2 concentration" ;
		CO2:units = "ppmv" ;
	float N2O(time) ;
		N2O:long_name = "Atmospheric N2O concentration" ;
		N2O:units = "ppbv" ;
	float year(time) ;
		year:long_name = "Year AD" ;

// global attributes:
		:description = "historical atmospheric CO2 and CH4 time series created on 2024/07/25/12:47:54; data source:Year:year,Value:number,Polutant:text\n" ;
data:

 CH4 = 712.7525, 712.8025, 714.8025, 717.9925, 717.1425, 713.7325, 712.0025, 
    715.6925, 724.6225, 728.6225, 727.7725, 730.1825, 712.9445, 712.9945, 
    714.9945, 718.1845, 717.3345, 713.9245, 712.1945, 715.8845, 724.8145, 
    728.8145, 727.9645, 730.3745, 713.1365, 713.1865, 715.1865, 718.3765, 
    717.5265, 714.1165, 712.3865, 716.0765, 725.0065, 729.0065, 728.1565, 
    730.5665, 713.3285, 713.3785, 715.3785, 718.5685, 717.7185, 714.3085, 
    712.5785, 716.2685, 725.1985, 729.1985, 728.3485, 730.7585, 713.5205, 
    713.5705, 715.5705, 718.7605, 717.9105, 714.5005, 712.7705, 716.4605, 
    725.3905, 729.3905, 728.5405, 730.9505, 713.7125, 713.7625, 715.7625, 
    718.9525, 718.1025, 714.6925, 712.9625, 716.6525, 725.5825, 729.5825, 
    728.7325, 731.1425, 713.9045, 713.9545, 715.9545, 719.1445, 718.2945, 
    714.8845, 713.1545, 716.8445, 725.7745, 729.7745, 728.9245, 731.3345, 
    714.0965, 714.1465, 716.1465, 719.3365, 718.4865, 715.0765, 713.3465, 
    717.0365, 725.9665, 729.9665, 729.1165, 731.5265, 714.2885, 714.3385, 
    716.3385, 719.5285, 718.6785, 715.2685, 713.5385, 717.2285, 726.1585, 
    730.1585, 729.3085, 731.7185, 714.4805, 714.5305, 716.5305, 719.7205, 
    718.8705, 715.4605, 713.7305, 717.4205, 726.3505, 730.3505, 729.5005, 
    731.9105, 714.6725, 714.7225, 716.7225, 719.9125, 719.0625, 715.6525, 
    713.9225, 717.6125, 726.5425, 730.5425, 729.6925, 732.1025, 715.2285, 
    715.2785, 717.2785, 720.4685, 719.6185, 716.2085, 714.4785, 718.1685, 
    727.0985, 731.0985, 730.2485, 732.6585, 715.7845, 715.8345, 717.8345, 
    721.0245, 720.1745, 716.7645, 715.0345, 718.7245, 727.6545, 731.6545, 
    730.8045, 733.2145, 716.3405, 716.3905, 718.3905, 721.5805, 720.7305, 
    717.3205, 715.5905, 719.2805, 728.2105, 732.2105, 731.3605, 733.7705, 
    716.8965, 716.9465, 718.9465, 722.1365, 721.2865, 717.8765, 716.1465, 
    719.8365, 728.7665, 732.7665, 731.9165, 734.3265, 717.4525, 717.5025, 
    719.5025, 722.6925, 721.8425, 718.4325, 716.7025, 720.3925, 729.3225, 
    733.3225, 732.4725, 734.8825, 718.0105, 718.0605, 720.0605, 723.2505, 
    722.4005, 718.9905, 717.2605, 720.9505, 729.8805, 733.8805, 733.0305, 
    735.4405, 718.5685, 718.6185, 720.6185, 723.8085, 722.9585, 719.5485, 
    717.8185, 721.5085, 730.4385, 734.4385, 733.5885, 735.9985, 719.1265, 
    719.1765, 721.1765, 724.3665, 723.5165, 720.1065, 718.3765, 722.0665, 
    730.9965, 734.9965, 734.1465, 736.5565, 719.6845, 719.7345, 721.7345, 
    724.9245, 724.0745, 720.6645, 718.9345, 722.6245, 731.5545, 735.5545, 
    734.7045, 737.1145, 720.2425, 720.2925, 722.2925, 725.4825, 724.6325, 
    721.2225, 719.4925, 723.1825, 732.1125, 736.1125, 735.2625, 737.6725, 
    721.0485, 721.0985, 723.0985, 726.2885, 725.4385, 722.0285, 720.2985, 
    723.9885, 732.9185, 736.9185, 736.0685, 738.4785, 721.8545, 721.9045, 
    723.9045, 727.0945, 726.2445, 722.8345, 721.1045, 724.7945, 733.7245, 
    737.7245, 736.8745, 739.2845, 722.6605, 722.7105, 724.7105, 727.9005, 
    727.0505, 723.6405, 721.9105, 725.6005, 734.5305, 738.5305, 737.6805, 
    740.0905, 723.4665, 723.5165, 725.5165, 728.7065, 727.8565, 724.4465, 
    722.7165, 726.4065, 735.3365, 739.3365, 738.4865, 740.8965, 724.2725, 
    724.3225, 726.3225, 729.5125, 728.6625, 725.2525, 723.5225, 727.2125, 
    736.1425, 740.1425, 739.2925, 741.7025, 725.0805, 725.1305, 727.1305, 
    730.3205, 729.4705, 726.0605, 724.3305, 728.0205, 736.9505, 740.9505, 
    740.1005, 742.5105, 725.8885, 725.9385, 727.9385, 731.1285, 730.2785, 
    726.8685, 725.1385, 728.8285, 737.7585, 741.7585, 740.9085, 743.3185, 
    726.6965, 726.7465, 728.7465, 731.9365, 731.0865, 727.6765, 725.9465, 
    729.6365, 738.5665, 742.5665, 741.7165, 744.1265, 727.5045, 727.5545, 
    729.5545, 732.7445, 731.8945, 728.4845, 726.7545, 730.4445, 739.3745, 
    743.3745, 742.5245, 744.9345, 728.3125, 728.3625, 730.3625, 733.5525, 
    732.7025, 729.2925, 727.5625, 731.2525, 740.1825, 744.1825, 743.3325, 
    745.7425, 729.2565, 729.3065, 731.3065, 734.4965, 733.6465, 730.2365, 
    728.5065, 732.1965, 741.1265, 745.1265, 744.2765, 746.6865, 730.2005, 
    730.2505, 732.2505, 735.4405, 734.5905, 731.1805, 729.4505, 733.1405, 
    742.0705, 746.0705, 745.2205, 747.6305, 731.1445, 731.1945, 733.1945, 
    736.3845, 735.5345, 732.1245, 730.3945, 734.0845, 743.0145, 747.0145, 
    746.1645, 748.5745, 732.0885, 732.1385, 734.1385, 737.3285, 736.4785, 
    733.0685, 731.3385, 735.0285, 743.9585, 747.9585, 747.1085, 749.5185, 
    733.0325, 733.0825, 735.0825, 738.2725, 737.4225, 734.0125, 732.2825, 
    735.9725, 744.9025, 748.9025, 748.0525, 750.4625, 733.9765, 734.0265, 
    736.0265, 739.2165, 738.3665, 734.9565, 733.2265, 736.9165, 745.8465, 
    749.8465, 748.9965, 751.4065, 734.9205, 734.9705, 736.9705, 740.1605, 
    739.3105, 735.9005, 734.1705, 737.8605, 746.7905, 750.7905, 749.9405, 
    752.3505, 735.8645, 735.9145, 737.9145, 741.1045, 740.2545, 736.8445, 
    735.1145, 738.8045, 747.7345, 751.7345, 750.8845, 753.2945, 736.8085, 
    736.8585, 738.8585, 742.0485, 741.1985, 737.7885, 736.0585, 739.7485, 
    748.6785, 752.6785, 751.8285, 754.2385, 737.7525, 737.8025, 739.8025, 
    742.9925, 742.1425, 738.7325, 737.0025, 740.6925, 749.6225, 753.6225, 
    752.7725, 755.1825, 738.4305, 738.4805, 740.4805, 743.6705, 742.8205, 
    739.4105, 737.6805, 741.3705, 750.3005, 754.3005, 753.4505, 755.8605, 
    739.1085, 739.1585, 741.1585, 744.3485, 743.4985, 740.0885, 738.3585, 
    742.0485, 750.9785, 754.9785, 754.1285, 756.5385, 739.7865, 739.8365, 
    741.8365, 745.0265, 744.1765, 740.7665, 739.0365, 742.7265, 751.6565, 
    755.6565, 754.8065, 757.2165, 740.4645, 740.5145, 742.5145, 745.7045, 
    744.8545, 741.4445, 739.7145, 743.4045, 752.3345, 756.3345, 755.4845, 
    757.8945, 741.1425, 741.1925, 743.1925, 746.3825, 745.5325, 742.1225, 
    740.3925, 744.0825, 753.0125, 757.0125, 756.1625, 758.5725, 741.8225, 
    741.8725, 743.8725, 747.0625, 746.2125, 742.8025, 741.0725, 744.7625, 
    753.6925, 757.6925, 756.8425, 759.2525, 742.5025, 742.5525, 744.5525, 
    747.7425, 746.8925, 743.4825, 741.7525, 745.4425, 754.3725, 758.3725, 
    757.5225, 759.9325, 743.1825, 743.2325, 745.2325, 748.4225, 747.5725, 
    744.1625, 742.4325, 746.1225, 755.0525, 759.0525, 758.2025, 760.6125, 
    743.8625, 743.9125, 745.9125, 749.1025, 748.2525, 744.8425, 743.1125, 
    746.8025, 755.7325, 759.7325, 758.8825, 761.2925, 744.5425, 744.5925, 
    746.5925, 749.7825, 748.9325, 745.5225, 743.7925, 747.4825, 756.4125, 
    760.4125, 759.5625, 761.9725, 745.4725, 745.5225, 747.5225, 750.7125, 
    749.8625, 746.4525, 744.7225, 748.4125, 757.3425, 761.3425, 760.4925, 
    762.9025, 746.4025, 746.4525, 748.4525, 751.6425, 750.7925, 747.3825, 
    745.6525, 749.3425, 758.2725, 762.2725, 761.4225, 763.8325, 747.3325, 
    747.3825, 749.3825, 752.5725, 751.7225, 748.3125, 746.5825, 750.2725, 
    759.2025, 763.2025, 762.3525, 764.7625, 748.2625, 748.3125, 750.3125, 
    753.5025, 752.6525, 749.2425, 747.5125, 751.2025, 760.1325, 764.1325, 
    763.2825, 765.6925, 749.1925, 749.2425, 751.2425, 754.4325, 753.5825, 
    750.1725, 748.4425, 752.1325, 761.0625, 765.0625, 764.2125, 766.6225, 
    750.1245, 750.1745, 752.1745, 755.3645, 754.5145, 751.1045, 749.3745, 
    753.0645, 761.9945, 765.9945, 765.1445, 767.5545, 751.0565, 751.1065, 
    753.1065, 756.2965, 755.4465, 752.0365, 750.3065, 753.9965, 762.9265, 
    766.9265, 766.0765, 768.4865, 751.9885, 752.0385, 754.0385, 757.2285, 
    756.3785, 752.9685, 751.2385, 754.9285, 763.8585, 767.8585, 767.0085, 
    769.4185, 752.9205, 752.9705, 754.9705, 758.1605, 757.3105, 753.9005, 
    752.1705, 755.8605, 764.7905, 768.7905, 767.9405, 770.3505, 753.8525, 
    753.9025, 755.9025, 759.0925, 758.2425, 754.8325, 753.1025, 756.7925, 
    765.7225, 769.7225, 768.8725, 771.2825, 754.8145, 754.8645, 756.8645, 
    760.0545, 759.2045, 755.7945, 754.0645, 757.7545, 766.6845, 770.6845, 
    769.8345, 772.2445, 755.7765, 755.8265, 757.8265, 761.0165, 760.1665, 
    756.7565, 755.0265, 758.7165, 767.6465, 771.6465, 770.7965, 773.2065, 
    756.7385, 756.7885, 758.7885, 761.9785, 761.1285, 757.7185, 755.9885, 
    759.6785, 768.6085, 772.6085, 771.7585, 774.1685, 757.7005, 757.7505, 
    759.7505, 762.9405, 762.0905, 758.6805, 756.9505, 760.6405, 769.5705, 
    773.5705, 772.7205, 775.1305, 758.6625, 758.7125, 760.7125, 763.9025, 
    763.0525, 759.6425, 757.9125, 761.6025, 770.5325, 774.5325, 773.6825, 
    776.0925, 759.6245, 759.6745, 761.6745, 764.8645, 764.0145, 760.6045, 
    758.8745, 762.5645, 771.4945, 775.4945, 774.6445, 777.0545, 760.5865, 
    760.6365, 762.6365, 765.8265, 764.9765, 761.5665, 759.8365, 763.5265, 
    772.4565, 776.4565, 775.6065, 778.0165, 761.5485, 761.5985, 763.5985, 
    766.7885, 765.9385, 762.5285, 760.7985, 764.4885, 773.4185, 777.4185, 
    776.5685, 778.9785, 762.5105, 762.5605, 764.5605, 767.7505, 766.9005, 
    763.4905, 761.7605, 765.4505, 774.3805, 778.3805, 777.5305, 779.9405, 
    763.4725, 763.5225, 765.5225, 768.7125, 767.8625, 764.4525, 762.7225, 
    766.4125, 775.3425, 779.3425, 778.4925, 780.9025, 764.4345, 764.4845, 
    766.4845, 769.6745, 768.8245, 765.4145, 763.6845, 767.3745, 776.3045, 
    780.3045, 779.4545, 781.8645, 765.3965, 765.4465, 767.4465, 770.6365, 
    769.7865, 766.3765, 764.6465, 768.3365, 777.2665, 781.2665, 780.4165, 
    782.8265, 766.3585, 766.4085, 768.4085, 771.5985, 770.7485, 767.3385, 
    765.6085, 769.2985, 778.2285, 782.2285, 781.3785, 783.7885, 767.3205, 
    767.3705, 769.3705, 772.5605, 771.7105, 768.3005, 766.5705, 770.2605, 
    779.1905, 783.1905, 782.3405, 784.7505, 768.2825, 768.3325, 770.3325, 
    773.5225, 772.6725, 769.2625, 767.5325, 771.2225, 780.1525, 784.1525, 
    783.3025, 785.7125, 769.2445, 769.2945, 771.2945, 774.4845, 773.6345, 
    770.2245, 768.4945, 772.1845, 781.1145, 785.1145, 784.2645, 786.6745, 
    770.2065, 770.2565, 772.2565, 775.4465, 774.5965, 771.1865, 769.4565, 
    773.1465, 782.0765, 786.0765, 785.2265, 787.6365, 771.1685, 771.2185, 
    773.2185, 776.4085, 775.5585, 772.1485, 770.4185, 774.1085, 783.0385, 
    787.0385, 786.1885, 788.5985, 772.1305, 772.1805, 774.1805, 777.3705, 
    776.5205, 773.1105, 771.3805, 775.0705, 784.0005, 788.0005, 787.1505, 
    789.5605, 773.0925, 773.1425, 775.1425, 778.3325, 777.4825, 774.0725, 
    772.3425, 776.0325, 784.9625, 788.9625, 788.1125, 790.5225, 774.0645, 
    774.1145, 776.1145, 779.3045, 778.4545, 775.0445, 773.3145, 777.0045, 
    785.9345, 789.9345, 789.0845, 791.4945, 775.0365, 775.0865, 777.0865, 
    780.2765, 779.4265, 776.0165, 774.2865, 777.9765, 786.9065, 790.9065, 
    790.0565, 792.4665, 776.0085, 776.0585, 778.0585, 781.2485, 780.3985, 
    776.9885, 775.2585, 778.9485, 787.8785, 791.8785, 791.0285, 793.4385, 
    776.9805, 777.0305, 779.0305, 782.2205, 781.3705, 777.9605, 776.2305, 
    779.9205, 788.8505, 792.8505, 792.0005, 794.4105, 777.9525, 778.0025, 
    780.0025, 783.1925, 782.3425, 778.9325, 777.2025, 780.8925, 789.8225, 
    793.8225, 792.9725, 795.3825, 778.9225, 778.9725, 780.9725, 784.1625, 
    783.3125, 779.9025, 778.1725, 781.8625, 790.7925, 794.7925, 793.9425, 
    796.3525, 779.8925, 779.9425, 781.9425, 785.1325, 784.2825, 780.8725, 
    779.1425, 782.8325, 791.7625, 795.7625, 794.9125, 797.3225, 780.8625, 
    780.9125, 782.9125, 786.1025, 785.2525, 781.8425, 780.1125, 783.8025, 
    792.7325, 796.7325, 795.8825, 798.2925, 781.8325, 781.8825, 783.8825, 
    787.0725, 786.2225, 782.8125, 781.0825, 784.7725, 793.7025, 797.7025, 
    796.8525, 799.2625, 782.8025, 782.8525, 784.8525, 788.0425, 787.1925, 
    783.7825, 782.0525, 785.7425, 794.6725, 798.6725, 797.8225, 800.2325, 
    784.0385, 784.0885, 786.0885, 789.2785, 788.4285, 785.0185, 783.2885, 
    786.9785, 795.9085, 799.9085, 799.0585, 801.4685, 785.2745, 785.3245, 
    787.3245, 790.5145, 789.6645, 786.2545, 784.5245, 788.2145, 797.1445, 
    801.1445, 800.2945, 802.7045, 786.5105, 786.5605, 788.5605, 791.7505, 
    790.9005, 787.4905, 785.7605, 789.4505, 798.3805, 802.3805, 801.5305, 
    803.9405, 787.7465, 787.7965, 789.7965, 792.9865, 792.1365, 788.7265, 
    786.9965, 790.6865, 799.6165, 803.6165, 802.7665, 805.1765, 788.9825, 
    789.0325, 791.0325, 794.2225, 793.3725, 789.9625, 788.2325, 791.9225, 
    800.8525, 804.8525, 804.0025, 806.4125, 790.2185, 790.2685, 792.2685, 
    795.4585, 794.6085, 791.1985, 789.4685, 793.1585, 802.0885, 806.0885, 
    805.2385, 807.6485, 791.4545, 791.5045, 793.5045, 796.6945, 795.8445, 
    792.4345, 790.7045, 794.3945, 803.3245, 807.3245, 806.4745, 808.8845, 
    792.6905, 792.7405, 794.7405, 797.9305, 797.0805, 793.6705, 791.9405, 
    795.6305, 804.5605, 808.5605, 807.7105, 810.1205, 793.9265, 793.9765, 
    795.9765, 799.1665, 798.3165, 794.9065, 793.1765, 796.8665, 805.7965, 
    809.7965, 808.9465, 811.3565, 795.1625, 795.2125, 797.2125, 800.4025, 
    799.5525, 796.1425, 794.4125, 798.1025, 807.0325, 811.0325, 810.1825, 
    812.5925, 796.5785, 796.6285, 798.6285, 801.8185, 800.9685, 797.5585, 
    795.8285, 799.5185, 808.4485, 812.4485, 811.5985, 814.0085, 797.9945, 
    798.0445, 800.0445, 803.2345, 802.3845, 798.9745, 797.2445, 800.9345, 
    809.8645, 813.8645, 813.0145, 815.4245, 799.4105, 799.4605, 801.4605, 
    804.6505, 803.8005, 800.3905, 798.6605, 802.3505, 811.2805, 815.2805, 
    814.4305, 816.8405, 800.8265, 800.8765, 802.8765, 806.0665, 805.2165, 
    801.8065, 800.0765, 803.7665, 812.6965, 816.6965, 815.8465, 818.2565, 
    802.2425, 802.2925, 804.2925, 807.4825, 806.6325, 803.2225, 801.4925, 
    805.1825, 814.1125, 818.1125, 817.2625, 819.6725, 803.6605, 803.7105, 
    805.7105, 808.9005, 808.0505, 804.6405, 802.9105, 806.6005, 815.5305, 
    819.5305, 818.6805, 821.0905, 805.0785, 805.1285, 807.1285, 810.3185, 
    809.4685, 806.0585, 804.3285, 808.0185, 816.9485, 820.9485, 820.0985, 
    822.5085, 806.4965, 806.5465, 808.5465, 811.7365, 810.8865, 807.4765, 
    805.7465, 809.4365, 818.3665, 822.3665, 821.5165, 823.9265, 807.9145, 
    807.9645, 809.9645, 813.1545, 812.3045, 808.8945, 807.1645, 810.8545, 
    819.7845, 823.7845, 822.9345, 825.3445, 809.3325, 809.3825, 811.3825, 
    814.5725, 813.7225, 810.3125, 808.5825, 812.2725, 821.2025, 825.2025, 
    824.3525, 826.7625, 810.8905, 810.9405, 812.9405, 816.1305, 815.2805, 
    811.8705, 810.1405, 813.8305, 822.7605, 826.7605, 825.9105, 828.3205, 
    812.4485, 812.4985, 814.4985, 817.6885, 816.8385, 813.4285, 811.6985, 
    815.3885, 824.3185, 828.3185, 827.4685, 829.8785, 814.0065, 814.0565, 
    816.0565, 819.2465, 818.3965, 814.9865, 813.2565, 816.9465, 825.8765, 
    829.8765, 829.0265, 831.4365, 815.5645, 815.6145, 817.6145, 820.8045, 
    819.9545, 816.5445, 814.8145, 818.5045, 827.4345, 831.4345, 830.5845, 
    832.9945, 817.1225, 817.1725, 819.1725, 822.3625, 821.5125, 818.1025, 
    816.3725, 820.0625, 828.9925, 832.9925, 832.1425, 834.5525, 818.6825, 
    818.7325, 820.7325, 823.9225, 823.0725, 819.6625, 817.9325, 821.6225, 
    830.5525, 834.5525, 833.7025, 836.1125, 820.2425, 820.2925, 822.2925, 
    825.4825, 824.6325, 821.2225, 819.4925, 823.1825, 832.1125, 836.1125, 
    835.2625, 837.6725, 821.8025, 821.8525, 823.8525, 827.0425, 826.1925, 
    822.7825, 821.0525, 824.7425, 833.6725, 837.6725, 836.8225, 839.2325, 
    823.3625, 823.4125, 825.4125, 828.6025, 827.7525, 824.3425, 822.6125, 
    826.3025, 835.2325, 839.2325, 838.3825, 840.7925, 824.9225, 824.9725, 
    826.9725, 830.1625, 829.3125, 825.9025, 824.1725, 827.8625, 836.7925, 
    840.7925, 839.9425, 842.3525, 826.5525, 826.6025, 828.6025, 831.7925, 
    830.9425, 827.5325, 825.8025, 829.4925, 838.4225, 842.4225, 841.5725, 
    843.9825, 828.1825, 828.2325, 830.2325, 833.4225, 832.5725, 829.1625, 
    827.4325, 831.1225, 840.0525, 844.0525, 843.2025, 845.6125, 829.8125, 
    829.8625, 831.8625, 835.0525, 834.2025, 830.7925, 829.0625, 832.7525, 
    841.6825, 845.6825, 844.8325, 847.2425, 831.4425, 831.4925, 833.4925, 
    836.6825, 835.8325, 832.4225, 830.6925, 834.3825, 843.3125, 847.3125, 
    846.4625, 848.8725, 833.0725, 833.1225, 835.1225, 838.3125, 837.4625, 
    834.0525, 832.3225, 836.0125, 844.9425, 848.9425, 848.0925, 850.5025, 
    834.7025, 834.7525, 836.7525, 839.9425, 839.0925, 835.6825, 833.9525, 
    837.6425, 846.5725, 850.5725, 849.7225, 852.1325, 836.3325, 836.3825, 
    838.3825, 841.5725, 840.7225, 837.3125, 835.5825, 839.2725, 848.2025, 
    852.2025, 851.3525, 853.7625, 837.9625, 838.0125, 840.0125, 843.2025, 
    842.3525, 838.9425, 837.2125, 840.9025, 849.8325, 853.8325, 852.9825, 
    855.3925, 839.5925, 839.6425, 841.6425, 844.8325, 843.9825, 840.5725, 
    838.8425, 842.5325, 851.4625, 855.4625, 854.6125, 857.0225, 841.2225, 
    841.2725, 843.2725, 846.4625, 845.6125, 842.2025, 840.4725, 844.1625, 
    853.0925, 857.0925, 856.2425, 858.6525, 843.1965, 843.2465, 845.2465, 
    848.4365, 847.5865, 844.1765, 842.4465, 846.1365, 855.0665, 859.0665, 
    858.2165, 860.6265, 845.1705, 845.2205, 847.2205, 850.4105, 849.5605, 
    846.1505, 844.4205, 848.1105, 857.0405, 861.0405, 860.1905, 862.6005, 
    847.1445, 847.1945, 849.1945, 852.3845, 851.5345, 848.1245, 846.3945, 
    850.0845, 859.0145, 863.0145, 862.1645, 864.5745, 849.1185, 849.1685, 
    851.1685, 854.3585, 853.5085, 850.0985, 848.3685, 852.0585, 860.9885, 
    864.9885, 864.1385, 866.5485, 851.0925, 851.1425, 853.1425, 856.3325, 
    855.4825, 852.0725, 850.3425, 854.0325, 862.9625, 866.9625, 866.1125, 
    868.5225, 853.0665, 853.1165, 855.1165, 858.3065, 857.4565, 854.0465, 
    852.3165, 856.0065, 864.9365, 868.9365, 868.0865, 870.4965, 855.0405, 
    855.0905, 857.0905, 860.2805, 859.4305, 856.0205, 854.2905, 857.9805, 
    866.9105, 870.9105, 870.0605, 872.4705, 857.0145, 857.0645, 859.0645, 
    862.2545, 861.4045, 857.9945, 856.2645, 859.9545, 868.8845, 872.8845, 
    872.0345, 874.4445, 858.9885, 859.0385, 861.0385, 864.2285, 863.3785, 
    859.9685, 858.2385, 861.9285, 870.8585, 874.8585, 874.0085, 876.4185, 
    860.9625, 861.0125, 863.0125, 866.2025, 865.3525, 861.9425, 860.2125, 
    863.9025, 872.8325, 876.8325, 875.9825, 878.3925, 863.2705, 863.3205, 
    865.3205, 868.5105, 867.6605, 864.2505, 862.5205, 866.2105, 875.1405, 
    879.1405, 878.2905, 880.7005, 865.5785, 865.6285, 867.6285, 870.8185, 
    869.9685, 866.5585, 864.8285, 868.5185, 877.4485, 881.4485, 880.5985, 
    883.0085, 867.8865, 867.9365, 869.9365, 873.1265, 872.2765, 868.8665, 
    867.1365, 870.8265, 879.7565, 883.7565, 882.9065, 885.3165, 870.1945, 
    870.2445, 872.2445, 875.4345, 874.5845, 871.1745, 869.4445, 873.1345, 
    882.0645, 886.0645, 885.2145, 887.6245, 872.5025, 872.5525, 874.5525, 
    877.7425, 876.8925, 873.4825, 871.7525, 875.4425, 884.3725, 888.3725, 
    887.5225, 889.9325, 874.8105, 874.8605, 876.8605, 880.0505, 879.2005, 
    875.7905, 874.0605, 877.7505, 886.6805, 890.6805, 889.8305, 892.2405, 
    877.1185, 877.1685, 879.1685, 882.3585, 881.5085, 878.0985, 876.3685, 
    880.0585, 888.9885, 892.9885, 892.1385, 894.5485, 879.4265, 879.4765, 
    881.4765, 884.6665, 883.8165, 880.4065, 878.6765, 882.3665, 891.2965, 
    895.2965, 894.4465, 896.8565, 881.7345, 881.7845, 883.7845, 886.9745, 
    886.1245, 882.7145, 880.9845, 884.6745, 893.6045, 897.6045, 896.7545, 
    899.1645, 884.0425, 884.0925, 886.0925, 889.2825, 888.4325, 885.0225, 
    883.2925, 886.9825, 895.9125, 899.9125, 899.0625, 901.4725, 888.3965, 
    888.4465, 890.4465, 893.6365, 892.7865, 889.3765, 887.6465, 891.3365, 
    900.2665, 904.2665, 903.4165, 905.8265, 892.7505, 892.8005, 894.8005, 
    897.9905, 897.1405, 893.7305, 892.0005, 895.6905, 904.6205, 908.6205, 
    907.7705, 910.1805, 897.1045, 897.1545, 899.1545, 902.3445, 901.4945, 
    898.0845, 896.3545, 900.0445, 908.9745, 912.9745, 912.1245, 914.5345, 
    901.4585, 901.5085, 903.5085, 906.6985, 905.8485, 902.4385, 900.7085, 
    904.3985, 913.3285, 917.3285, 916.4785, 918.8885, 905.8125, 905.8625, 
    907.8625, 911.0525, 910.2025, 906.7925, 905.0625, 908.7525, 917.6825, 
    921.6825, 920.8325, 923.2425, 910.4905, 910.5405, 912.5405, 915.7305, 
    914.8805, 911.4705, 909.7405, 913.4305, 922.3605, 926.3605, 925.5105, 
    927.9205, 915.1685, 915.2185, 917.2185, 920.4085, 919.5585, 916.1485, 
    914.4185, 918.1085, 927.0385, 931.0385, 930.1885, 932.5985, 919.8465, 
    919.8965, 921.8965, 925.0865, 924.2365, 920.8265, 919.0965, 922.7865, 
    931.7165, 935.7165, 934.8665, 937.2765, 924.5245, 924.5745, 926.5745, 
    929.7645, 928.9145, 925.5045, 923.7745, 927.4645, 936.3945, 940.3945, 
    939.5445, 941.9545, 929.2025, 929.2525, 931.2525, 934.4425, 933.5925, 
    930.1825, 928.4525, 932.1425, 941.0725, 945.0725, 944.2225, 946.6325, 
    934.4065, 934.4565, 936.4565, 939.6465, 938.7965, 935.3865, 933.6565, 
    937.3465, 946.2765, 950.2765, 949.4265, 951.8365, 939.6105, 939.6605, 
    941.6605, 944.8505, 944.0005, 940.5905, 938.8605, 942.5505, 951.4805, 
    955.4805, 954.6305, 957.0405, 944.8145, 944.8645, 946.8645, 950.0545, 
    949.2045, 945.7945, 944.0645, 947.7545, 956.6845, 960.6845, 959.8345, 
    962.2445, 950.0185, 950.0685, 952.0685, 955.2585, 954.4085, 950.9985, 
    949.2685, 952.9585, 961.8885, 965.8885, 965.0385, 967.4485, 955.2225, 
    955.2725, 957.2725, 960.4625, 959.6125, 956.2025, 954.4725, 958.1625, 
    967.0925, 971.0925, 970.2425, 972.6525, 960.9725, 961.0225, 963.0225, 
    966.2125, 965.3625, 961.9525, 960.2225, 963.9125, 972.8425, 976.8425, 
    975.9925, 978.4025, 966.7225, 966.7725, 968.7725, 971.9625, 971.1125, 
    967.7025, 965.9725, 969.6625, 978.5925, 982.5925, 981.7425, 984.1525, 
    972.4725, 972.5225, 974.5225, 977.7125, 976.8625, 973.4525, 971.7225, 
    975.4125, 984.3425, 988.3425, 987.4925, 989.9025, 978.2225, 978.2725, 
    980.2725, 983.4625, 982.6125, 979.2025, 977.4725, 981.1625, 990.0925, 
    994.0925, 993.2425, 995.6525, 983.9725, 984.0225, 986.0225, 989.2125, 
    988.3625, 984.9525, 983.2225, 986.9125, 995.8425, 999.8425, 998.9925, 
    1001.403, 989.9665, 990.0165, 992.0165, 995.2065, 994.3565, 990.9465, 
    989.2165, 992.9065, 1001.836, 1005.836, 1004.987, 1007.396, 995.9605, 
    996.0105, 998.0105, 1001.201, 1000.351, 996.9405, 995.2105, 998.9005, 
    1007.831, 1011.831, 1010.981, 1013.391, 1001.955, 1002.005, 1004.005, 
    1007.195, 1006.344, 1002.935, 1001.205, 1004.894, 1013.825, 1017.825, 
    1016.974, 1019.385, 1007.948, 1007.998, 1009.998, 1013.188, 1012.339, 
    1008.929, 1007.198, 1010.888, 1019.818, 1023.818, 1022.969, 1025.379, 
    1013.943, 1013.992, 1015.992, 1019.182, 1018.333, 1014.922, 1013.193, 
    1016.883, 1025.812, 1029.812, 1028.963, 1031.373, 1019.713, 1019.763, 
    1021.763, 1024.953, 1024.103, 1020.693, 1018.963, 1022.653, 1031.583, 
    1035.583, 1034.733, 1037.142, 1025.483, 1025.532, 1027.532, 1030.723, 
    1029.873, 1026.463, 1024.733, 1028.422, 1037.353, 1041.353, 1040.502, 
    1042.912, 1031.252, 1031.302, 1033.302, 1036.493, 1035.642, 1032.233, 
    1030.502, 1034.193, 1043.123, 1047.123, 1046.272, 1048.682, 1037.022, 
    1037.073, 1039.073, 1042.262, 1041.412, 1038.002, 1036.272, 1039.963, 
    1048.892, 1052.892, 1052.042, 1054.453, 1042.792, 1042.843, 1044.843, 
    1048.032, 1047.182, 1043.772, 1042.042, 1045.733, 1054.662, 1058.662, 
    1057.812, 1060.223, 1048.291, 1048.34, 1050.34, 1053.531, 1052.681, 
    1049.271, 1047.541, 1051.23, 1060.161, 1064.161, 1063.311, 1065.72, 
    1053.788, 1053.839, 1055.839, 1059.028, 1058.178, 1054.769, 1053.038, 
    1056.729, 1065.658, 1069.658, 1068.808, 1071.219, 1059.286, 1059.337, 
    1061.337, 1064.526, 1063.677, 1060.266, 1058.536, 1062.226, 1071.156, 
    1075.156, 1074.307, 1076.717, 1064.785, 1064.834, 1066.834, 1070.025, 
    1069.175, 1065.765, 1064.035, 1067.724, 1076.655, 1080.655, 1079.804, 
    1082.214, 1070.282, 1070.333, 1072.333, 1075.522, 1074.672, 1071.262, 
    1069.532, 1073.223, 1082.152, 1086.152, 1085.302, 1087.713, 1075.454, 
    1075.505, 1077.505, 1080.694, 1079.844, 1076.434, 1074.704, 1078.395, 
    1087.324, 1091.324, 1090.474, 1092.885, 1080.626, 1080.677, 1082.677, 
    1085.866, 1085.016, 1081.606, 1079.876, 1083.567, 1092.496, 1096.496, 
    1095.646, 1098.057, 1085.798, 1085.849, 1087.849, 1091.038, 1090.188, 
    1086.778, 1085.048, 1088.739, 1097.668, 1101.668, 1100.818, 1103.229, 
    1090.97, 1091.021, 1093.021, 1096.21, 1095.36, 1091.95, 1090.22, 
    1093.911, 1102.84, 1106.84, 1105.99, 1108.401, 1096.142, 1096.193, 
    1098.193, 1101.382, 1100.532, 1097.123, 1095.392, 1099.083, 1108.012, 
    1112.012, 1111.162, 1113.573, 1101.428, 1101.479, 1103.479, 1106.668, 
    1105.818, 1102.408, 1100.678, 1104.369, 1113.298, 1117.298, 1116.448, 
    1118.859, 1106.714, 1106.765, 1108.765, 1111.954, 1111.104, 1107.694, 
    1105.964, 1109.655, 1118.584, 1122.584, 1121.734, 1124.145, 1112, 
    1112.051, 1114.051, 1117.24, 1116.391, 1112.98, 1111.25, 1114.941, 
    1123.87, 1127.87, 1127.021, 1129.431, 1117.286, 1117.337, 1119.337, 
    1122.526, 1121.677, 1118.266, 1116.536, 1120.226, 1129.156, 1133.156, 
    1132.307, 1134.717, 1122.573, 1122.623, 1124.623, 1127.812, 1126.963, 
    1123.552, 1121.823, 1125.512, 1134.443, 1138.443, 1137.593, 1140.002, 
    1129.152, 1129.203, 1131.203, 1134.392, 1133.542, 1130.132, 1128.402, 
    1132.093, 1141.022, 1145.022, 1144.172, 1146.583, 1135.733, 1135.782, 
    1137.782, 1140.973, 1140.123, 1136.713, 1134.983, 1138.672, 1147.603, 
    1151.603, 1150.752, 1153.162, 1142.312, 1142.363, 1144.363, 1147.552, 
    1146.703, 1143.292, 1141.562, 1145.252, 1154.182, 1158.182, 1157.333, 
    1159.743, 1148.892, 1148.943, 1150.943, 1154.132, 1153.282, 1149.873, 
    1148.142, 1151.833, 1160.762, 1164.762, 1163.912, 1166.323, 1155.473, 
    1155.522, 1157.522, 1160.713, 1159.863, 1156.453, 1154.723, 1158.412, 
    1167.343, 1171.343, 1170.493, 1172.902, 1164.532, 1164.583, 1166.583, 
    1169.772, 1168.922, 1165.512, 1163.782, 1167.473, 1176.402, 1180.402, 
    1179.552, 1181.963, 1173.593, 1173.642, 1175.642, 1178.833, 1177.983, 
    1174.573, 1172.843, 1176.532, 1185.463, 1189.463, 1188.613, 1191.022, 
    1182.652, 1182.703, 1184.703, 1187.892, 1187.042, 1183.632, 1181.902, 
    1185.593, 1194.522, 1198.522, 1197.672, 1200.083, 1191.713, 1191.762, 
    1193.762, 1196.953, 1196.103, 1192.693, 1190.963, 1194.652, 1203.583, 
    1207.583, 1206.733, 1209.142, 1200.772, 1200.823, 1202.823, 1206.012, 
    1205.162, 1201.752, 1200.022, 1203.713, 1212.642, 1216.642, 1215.792, 
    1218.203, 1211.96, 1212.01, 1214.01, 1217.2, 1216.35, 1212.941, 1211.21, 
    1214.901, 1223.83, 1227.83, 1226.98, 1229.391, 1223.149, 1223.198, 
    1225.198, 1228.389, 1227.538, 1224.129, 1222.399, 1226.089, 1235.019, 
    1239.019, 1238.168, 1240.578, 1234.337, 1234.386, 1236.386, 1239.577, 
    1238.726, 1235.317, 1233.587, 1237.276, 1246.207, 1250.207, 1249.356, 
    1251.766, 1245.525, 1245.574, 1247.574, 1250.765, 1249.915, 1246.505, 
    1244.775, 1248.464, 1257.395, 1261.395, 1260.545, 1262.954, 1256.713, 
    1256.762, 1258.762, 1261.953, 1261.103, 1257.693, 1255.963, 1259.652, 
    1268.583, 1272.583, 1271.733, 1274.142, 1269.812, 1269.863, 1271.863, 
    1275.052, 1274.203, 1270.792, 1269.062, 1272.752, 1281.682, 1285.682, 
    1284.833, 1287.243, 1282.912, 1282.963, 1284.963, 1288.152, 1287.302, 
    1283.892, 1282.162, 1285.853, 1294.782, 1298.782, 1297.932, 1300.343, 
    1296.012, 1296.062, 1298.062, 1301.252, 1300.402, 1296.993, 1295.262, 
    1298.953, 1307.882, 1311.882, 1311.032, 1313.443, 1309.113, 1309.162, 
    1311.162, 1314.353, 1313.502, 1310.093, 1308.363, 1312.052, 1320.983, 
    1324.983, 1324.132, 1326.542, 1322.213, 1322.262, 1324.262, 1327.453, 
    1326.603, 1323.193, 1321.463, 1325.152, 1334.083, 1338.083, 1337.233, 
    1339.642, 1337.156, 1337.207, 1339.207, 1342.396, 1341.547, 1338.136, 
    1336.406, 1340.097, 1349.026, 1353.026, 1352.177, 1354.587, 1352.1, 
    1352.151, 1354.151, 1357.34, 1356.49, 1353.08, 1351.35, 1355.041, 
    1363.97, 1367.97, 1367.12, 1369.531, 1367.045, 1367.094, 1369.094, 
    1372.285, 1371.434, 1368.025, 1366.295, 1369.984, 1378.915, 1382.915, 
    1382.064, 1384.474, 1381.989, 1382.038, 1384.038, 1387.229, 1386.379, 
    1382.969, 1381.239, 1384.928, 1393.859, 1397.859, 1397.009, 1399.418, 
    1396.932, 1396.983, 1398.983, 1402.172, 1401.323, 1397.912, 1396.182, 
    1399.873, 1408.802, 1412.802, 1411.953, 1414.363, 1413.009, 1413.058, 
    1415.058, 1418.249, 1417.399, 1413.989, 1412.259, 1415.948, 1424.879, 
    1428.879, 1428.028, 1430.438, 1429.084, 1429.135, 1431.135, 1434.324, 
    1433.474, 1430.064, 1428.334, 1432.025, 1440.954, 1444.954, 1444.104, 
    1446.515, 1445.161, 1445.21, 1447.21, 1450.401, 1449.551, 1446.141, 
    1444.411, 1448.1, 1457.031, 1461.031, 1460.181, 1462.59, 1461.236, 
    1461.286, 1463.286, 1466.476, 1465.626, 1462.217, 1460.486, 1464.177, 
    1473.106, 1477.106, 1476.256, 1478.667, 1477.312, 1477.363, 1479.363, 
    1482.552, 1481.703, 1478.292, 1476.562, 1480.252, 1489.182, 1493.182, 
    1492.333, 1494.743, 1493.713, 1493.762, 1495.762, 1498.953, 1498.103, 
    1494.693, 1492.963, 1496.652, 1505.583, 1509.583, 1508.733, 1511.142, 
    1510.113, 1510.162, 1512.162, 1515.353, 1514.502, 1511.093, 1509.363, 
    1513.052, 1521.983, 1525.983, 1525.132, 1527.542, 1526.512, 1526.562, 
    1528.562, 1531.752, 1530.902, 1527.493, 1525.762, 1529.453, 1538.382, 
    1542.382, 1541.532, 1543.943, 1543.272, 1543.323, 1545.323, 1548.512, 
    1547.662, 1544.252, 1542.522, 1546.213, 1555.142, 1559.142, 1558.292, 
    1560.703, 1560.022, 1560.073, 1562.073, 1565.262, 1564.412, 1561.002, 
    1559.272, 1562.963, 1571.892, 1575.892, 1575.042, 1577.453, 1577.223, 
    1577.272, 1579.272, 1582.463, 1581.613, 1578.203, 1576.473, 1580.162, 
    1589.093, 1593.093, 1592.243, 1594.652, 1594.432, 1594.483, 1596.483, 
    1599.672, 1598.823, 1595.412, 1593.682, 1597.373, 1606.302, 1610.302, 
    1609.453, 1611.863, 1611.632, 1611.682, 1613.682, 1616.873, 1616.022, 
    1612.613, 1610.882, 1614.573, 1623.502, 1627.502, 1626.652, 1629.062, 
    1638.432, 1638.483, 1640.483, 1643.672, 1642.823, 1639.412, 1637.682, 
    1641.373, 1650.302, 1654.302, 1653.453, 1655.863, 1655.521, 1652.141, 
    1654.501, 1658.121, 1655.781, 1649.951, 1646.731, 1652.151, 1662.391, 
    1667.421, 1666.701, 1665.951, 1666.168, 1666.778, 1669.118, 1670.688, 
    1668.308, 1664.628, 1662.208, 1664.238, 1672.448, 1678.558, 1678.838, 
    1678.978, 1679.335, 1678.935, 1679.925, 1681.275, 1681.755, 1679.895, 
    1675.885, 1677.055, 1685.505, 1691.505, 1691.055, 1690.395, 1691.955, 
    1692.465, 1691.235, 1689.985, 1688.965, 1687.025, 1685.885, 1689.285, 
    1695.985, 1701.015, 1702.695, 1701.785, 1700.479, 1700.979, 1702.369, 
    1703.519, 1703.279, 1700.119, 1698.129, 1701.889, 1707.099, 1710.449, 
    1713.019, 1713.149, 1712.015, 1713.365, 1714.245, 1712.425, 1710.485, 
    1708.305, 1706.415, 1710.055, 1717.435, 1721.865, 1723.295, 1723.135, 
    1721.576, 1721.206, 1722.016, 1722.376, 1722.046, 1718.846, 1715.946, 
    1719.086, 1726.026, 1732.696, 1737.426, 1739.556, 1738.973, 1737.403, 
    1736.943, 1736.713, 1735.013, 1731.603, 1728.863, 1730.363, 1734.653, 
    1737.723, 1739.263, 1738.603, 1735.75, 1734.3, 1735.32, 1736.56, 1734.94, 
    1730.82, 1727.98, 1731.08, 1738.4, 1743.34, 1745.15, 1744.24, 1741.37, 
    1740.79, 1741.86, 1741.88, 1740.55, 1736.8, 1732.33, 1733.98, 1742.81, 
    1749.69, 1751.13, 1751.53, 1751.064, 1749.394, 1748.894, 1749.354, 
    1747.554, 1742.734, 1740.084, 1743.494, 1749.694, 1754.274, 1755.404, 
    1753.774, 1752.379, 1752.859, 1752.359, 1749.739, 1748.429, 1746.169, 
    1742.189, 1744.409, 1752.759, 1759.029, 1760.149, 1757.049, 1753.367, 
    1753.797, 1755.617, 1755.507, 1753.757, 1750.037, 1746.017, 1747.697, 
    1754.927, 1760.257, 1761.657, 1761.847, 1761.345, 1761.315, 1762.815, 
    1764.605, 1764.125, 1760.205, 1756.055, 1760.075, 1770.545, 1776.125, 
    1775.345, 1773.925, 1773.853, 1773.922, 1774.613, 1775.022, 1772.693, 
    1767.373, 1763.002, 1764.652, 1771.042, 1776.662, 1778.573, 1777.272, 
    1775.696, 1775.596, 1776.636, 1777.396, 1774.726, 1768.286, 1763.646, 
    1765.616, 1772.206, 1777.276, 1777.886, 1775.476, 1772.892, 1772.502, 
    1773.642, 1773.882, 1770.743, 1765.833, 1762.782, 1764.292, 1770.353, 
    1775.493, 1776.552, 1775.912, 1774.107, 1772.797, 1773.377, 1772.757, 
    1770.287, 1766.887, 1764.217, 1766.837, 1773.647, 1778.257, 1779.477, 
    1779.637, 1777.526, 1774.776, 1774.806, 1775.786, 1774.416, 1771.646, 
    1770.686, 1774.256, 1780.526, 1784.666, 1785.226, 1783.526, 1780.902, 
    1779.963, 1780.963, 1780.743, 1777.583, 1772.302, 1768.062, 1769.792, 
    1775.512, 1779.713, 1780.483, 1778.343, 1776.04, 1775.57, 1775.42, 
    1774.66, 1772.35, 1768.65, 1766.27, 1768, 1773.09, 1778.44, 1781.08, 
    1780.11, 1779.525, 1779.435, 1777.365, 1776.115, 1774.895, 1769.205, 
    1764.165, 1767.215, 1774.575, 1778.235, 1779.005, 1779.905, 1779.162, 
    1778.522, 1780.162, 1781.062, 1779.402, 1775.542, 1772.532, 1777.123, 
    1785.802, 1789.792, 1789.453, 1788.123, 1786.615, 1785.705, 1786.055, 
    1786.815, 1785.115, 1780.375, 1777.575, 1780.965, 1787.575, 1793.605, 
    1797.205, 1796.515, 1795.073, 1795.552, 1795.902, 1795.542, 1792.363, 
    1786.912, 1785.012, 1788.873, 1794.792, 1797.993, 1797.823, 1796.642, 
    1797.061, 1798.681, 1799.361, 1799.521, 1797.541, 1792.381, 1789.361, 
    1794.011, 1801.781, 1806.521, 1806.951, 1803.511, 1800.393, 1800.073, 
    1800.873, 1802.833, 1803.233, 1799.063, 1796.153, 1798.993, 1803.983, 
    1809.493, 1812.273, 1809.953, 1807.241, 1808.201, 1809.881, 1808.341, 
    1804.601, 1800.841, 1799.231, 1803.141, 1809.991, 1814.691, 1815.781, 
    1814.421, 1813.998, 1814.047, 1813.157, 1812.757, 1811.848, 1808.517, 
    1805.917, 1808.448, 1814.167, 1818.438, 1820.248, 1819.257, 1816.778, 
    1816.248, 1818.008, 1820.828, 1821.818, 1818.228, 1815.478, 1819.628, 
    1826.748, 1831.138, 1832.938, 1833.478, 1833.043, 1832.843, 1833.133, 
    1833.133, 1831.473, 1827.063, 1824.543, 1828.923, 1836.173, 1841.443, 
    1844.523, 1844.703, 1842.393, 1841.603, 1842.943, 1843.733, 1842.093, 
    1837.793, 1834.153, 1836.663, 1844.153, 1849.853, 1851.393, 1851.023, 
    1849.747, 1848.417, 1848.207, 1848.597, 1847.177, 1842.967, 1840.437, 
    1844.647, 1852.737, 1858.027, 1858.537, 1856.547, 1854.327, 1854.827, 
    1856.717, 1856.567, 1854.677, 1851.867, 1848.967, 1851.787, 1860.347, 
    1865.637, 1866.117, 1865.887, 1864.929, 1864.939, 1866.229, 1865.259, 
    1861.899, 1858.709, 1858.179, 1862.829, 1870.709, 1875.329, 1875.469, 
    1874.599, 1873.007, 1872.578, 1874.557, 1875.738, 1874.157, 1871.698, 
    1871.358, 1876.377, 1884.517, 1889.958, 1891.738, 1891.718, 1889.554, 
    1887.454, 1888.504, 1891.094, 1891.424, 1888.184, 1886.164, 1892.464, 
    1902.504, 1907.994, 1909.514, 1908.624, 1907.348, 1907.518, 1908.708, 
    1909.398, 1907.718, 1905.038, 1904.338, 1908.648, 1915.368, 1920.018, 
    1923.578, 1924.398, 1922.440, 1920.350, 1919.700, 1920.550, 1919.750,
    1915.650, 1913.990, 1917.990, 1925.310, 1930.570, 1931.780, 1931.880 ;

 CO2 = 277.7092, 278.4392, 279.0292, 279.4692, 279.4092, 278.5292, 276.7092, 
    275.5192, 276.1692, 277.5092, 278.5092, 278.9992, 277.7092, 278.4392, 
    279.0292, 279.4692, 279.4092, 278.5292, 276.7092, 275.5192, 276.1692, 
    277.5092, 278.5092, 278.9992, 277.7092, 278.4392, 279.0292, 279.4692, 
    279.4092, 278.5292, 276.7092, 275.5192, 276.1692, 277.5092, 278.5092, 
    278.9992, 277.7092, 278.4392, 279.0292, 279.4692, 279.4092, 278.5292, 
    276.7092, 275.5192, 276.1692, 277.5092, 278.5092, 278.9992, 277.7092, 
    278.4392, 279.0292, 279.4692, 279.4092, 278.5292, 276.7092, 275.5192, 
    276.1692, 277.5092, 278.5092, 278.9992, 277.7092, 278.4392, 279.0292, 
    279.4692, 279.4092, 278.5292, 276.7092, 275.5192, 276.1692, 277.5092, 
    278.5092, 278.9992, 277.7092, 278.4392, 279.0292, 279.4692, 279.4092, 
    278.5292, 276.7092, 275.5192, 276.1692, 277.5092, 278.5092, 278.9992, 
    277.7092, 278.4392, 279.0292, 279.4692, 279.4092, 278.5292, 276.7092, 
    275.5192, 276.1692, 277.5092, 278.5092, 278.9992, 277.7092, 278.4392, 
    279.0292, 279.4692, 279.4092, 278.5292, 276.7092, 275.5192, 276.1692, 
    277.5092, 278.5092, 278.9992, 277.7092, 278.4392, 279.0292, 279.4692, 
    279.4092, 278.5292, 276.7092, 275.5192, 276.1692, 277.5092, 278.5092, 
    278.9992, 277.7092, 278.4392, 279.0292, 279.4692, 279.4092, 278.5292, 
    276.7092, 275.5192, 276.1692, 277.5092, 278.5092, 278.9992, 277.7092, 
    278.4392, 279.0292, 279.4692, 279.4092, 278.5292, 276.7092, 275.5192, 
    276.1692, 277.5092, 278.5092, 278.9992, 277.7092, 278.4392, 279.0292, 
    279.4692, 279.4092, 278.5292, 276.7092, 275.5192, 276.1692, 277.5092, 
    278.5092, 278.9992, 277.7092, 278.4392, 279.0292, 279.4692, 279.4092, 
    278.5292, 276.7092, 275.5192, 276.1692, 277.5092, 278.5092, 278.9992, 
    277.7092, 278.4392, 279.0292, 279.4692, 279.4092, 278.5292, 276.7092, 
    275.5192, 276.1692, 277.5092, 278.5092, 278.9992, 277.7092, 278.4392, 
    279.0292, 279.4692, 279.4092, 278.5292, 276.7092, 275.5192, 276.1692, 
    277.5092, 278.5092, 278.9992, 277.8292, 278.5592, 279.1492, 279.5892, 
    279.5292, 278.6492, 276.8292, 275.6392, 276.2892, 277.6292, 278.6292, 
    279.1192, 277.9492, 278.6792, 279.2692, 279.7092, 279.6492, 278.7692, 
    276.9492, 275.7592, 276.4092, 277.7492, 278.7492, 279.2392, 278.0692, 
    278.7992, 279.3892, 279.8292, 279.7692, 278.8892, 277.0692, 275.8792, 
    276.5292, 277.8692, 278.8692, 279.3592, 278.1892, 278.9192, 279.5092, 
    279.9492, 279.8892, 279.0092, 277.1892, 275.9992, 276.6492, 277.9892, 
    278.9892, 279.4792, 278.3092, 279.0392, 279.6292, 280.0692, 280.0092, 
    279.1292, 277.3092, 276.1192, 276.7692, 278.1092, 279.1092, 279.5992, 
    278.4492, 279.1792, 279.7692, 280.2092, 280.1492, 279.2692, 277.4492, 
    276.2592, 276.9092, 278.2492, 279.2492, 279.7392, 278.5892, 279.3192, 
    279.9092, 280.3492, 280.2892, 279.4092, 277.5892, 276.3992, 277.0492, 
    278.3892, 279.3892, 279.8792, 278.7292, 279.4592, 280.0492, 280.4892, 
    280.4292, 279.5492, 277.7292, 276.5392, 277.1892, 278.5292, 279.5292, 
    280.0192, 278.8692, 279.5992, 280.1892, 280.6292, 280.5692, 279.6892, 
    277.8692, 276.6792, 277.3292, 278.6692, 279.6692, 280.1592, 279.0092, 
    279.7392, 280.3292, 280.7692, 280.7092, 279.8292, 278.0092, 276.8192, 
    277.4692, 278.8092, 279.8092, 280.2992, 279.1692, 279.8992, 280.4892, 
    280.9292, 280.8692, 279.9892, 278.1692, 276.9792, 277.6292, 278.9692, 
    279.9692, 280.4592, 279.3292, 280.0592, 280.6492, 281.0892, 281.0292, 
    280.1492, 278.3292, 277.1392, 277.7892, 279.1292, 280.1292, 280.6192, 
    279.4892, 280.2192, 280.8092, 281.2492, 281.1892, 280.3092, 278.4892, 
    277.2992, 277.9492, 279.2892, 280.2892, 280.7792, 279.6492, 280.3792, 
    280.9692, 281.4092, 281.3492, 280.4692, 278.6492, 277.4592, 278.1092, 
    279.4492, 280.4492, 280.9392, 279.8092, 280.5392, 281.1292, 281.5692, 
    281.5092, 280.6292, 278.8092, 277.6192, 278.2692, 279.6092, 280.6092, 
    281.0992, 279.9492, 280.6792, 281.2692, 281.7092, 281.6492, 280.7692, 
    278.9492, 277.7592, 278.4092, 279.7492, 280.7492, 281.2392, 280.0892, 
    280.8192, 281.4092, 281.8492, 281.7892, 280.9092, 279.0892, 277.8992, 
    278.5492, 279.8892, 280.8892, 281.3792, 280.2292, 280.9592, 281.5492, 
    281.9892, 281.9292, 281.0492, 279.2292, 278.0392, 278.6892, 280.0292, 
    281.0292, 281.5192, 280.3692, 281.0992, 281.6892, 282.1292, 282.0692, 
    281.1892, 279.3692, 278.1792, 278.8292, 280.1692, 281.1692, 281.6592, 
    280.5092, 281.2392, 281.8292, 282.2692, 282.2092, 281.3292, 279.5092, 
    278.3192, 278.9692, 280.3092, 281.3092, 281.7992, 280.6692, 281.3992, 
    281.9892, 282.4292, 282.3692, 281.4892, 279.6692, 278.4792, 279.1292, 
    280.4692, 281.4692, 281.9592, 280.8292, 281.5592, 282.1492, 282.5892, 
    282.5292, 281.6492, 279.8292, 278.6392, 279.2892, 280.6292, 281.6292, 
    282.1192, 280.9892, 281.7192, 282.3092, 282.7492, 282.6892, 281.8092, 
    279.9892, 278.7992, 279.4492, 280.7892, 281.7892, 282.2792, 281.1492, 
    281.8792, 282.4692, 282.9092, 282.8492, 281.9692, 280.1492, 278.9592, 
    279.6092, 280.9492, 281.9492, 282.4392, 281.3092, 282.0392, 282.6292, 
    283.0692, 283.0092, 282.1292, 280.3092, 279.1192, 279.7692, 281.1092, 
    282.1092, 282.5992, 281.4492, 282.1792, 282.7692, 283.2092, 283.1492, 
    282.2692, 280.4492, 279.2592, 279.9092, 281.2492, 282.2492, 282.7392, 
    281.5892, 282.3192, 282.9092, 283.3492, 283.2892, 282.4092, 280.5892, 
    279.3992, 280.0492, 281.3892, 282.3892, 282.8792, 281.7292, 282.4592, 
    283.0492, 283.4892, 283.4292, 282.5492, 280.7292, 279.5392, 280.1892, 
    281.5292, 282.5292, 283.0192, 281.8692, 282.5992, 283.1892, 283.6292, 
    283.5692, 282.6892, 280.8692, 279.6792, 280.3292, 281.6692, 282.6692, 
    283.1592, 282.0092, 282.7392, 283.3292, 283.7692, 283.7092, 282.8292, 
    281.0092, 279.8192, 280.4692, 281.8092, 282.8092, 283.2992, 282.1292, 
    282.8592, 283.4492, 283.8892, 283.8292, 282.9492, 281.1292, 279.9392, 
    280.5892, 281.9292, 282.9292, 283.4192, 282.2492, 282.9792, 283.5692, 
    284.0092, 283.9492, 283.0692, 281.2492, 280.0592, 280.7092, 282.0492, 
    283.0492, 283.5392, 282.3692, 283.0992, 283.6892, 284.1292, 284.0692, 
    283.1892, 281.3692, 280.1792, 280.8292, 282.1692, 283.1692, 283.6592, 
    282.4892, 283.2192, 283.8092, 284.2492, 284.1892, 283.3092, 281.4892, 
    280.2992, 280.9492, 282.2892, 283.2892, 283.7792, 282.6092, 283.3392, 
    283.9292, 284.3692, 284.3092, 283.4292, 281.6092, 280.4192, 281.0692, 
    282.4092, 283.4092, 283.8992, 282.7092, 283.4392, 284.0292, 284.4692, 
    284.4092, 283.5292, 281.7092, 280.5192, 281.1692, 282.5092, 283.5092, 
    283.9992, 282.8092, 283.5392, 284.1292, 284.5692, 284.5092, 283.6292, 
    281.8092, 280.6192, 281.2692, 282.6092, 283.6092, 284.0992, 282.9092, 
    283.6392, 284.2292, 284.6692, 284.6092, 283.7292, 281.9092, 280.7192, 
    281.3692, 282.7092, 283.7092, 284.1992, 283.0092, 283.7392, 284.3292, 
    284.7692, 284.7092, 283.8292, 282.0092, 280.8192, 281.4692, 282.8092, 
    283.8092, 284.2992, 283.1092, 283.8392, 284.4292, 284.8692, 284.8092, 
    283.9292, 282.1092, 280.9192, 281.5692, 282.9092, 283.9092, 284.3992, 
    283.1892, 283.9192, 284.5092, 284.9492, 284.8892, 284.0092, 282.1892, 
    280.9992, 281.6492, 282.9892, 283.9892, 284.4792, 283.2692, 283.9992, 
    284.5892, 285.0292, 284.9692, 284.0892, 282.2692, 281.0792, 281.7292, 
    283.0692, 284.0692, 284.5592, 283.3492, 284.0792, 284.6692, 285.1092, 
    285.0492, 284.1692, 282.3492, 281.1592, 281.8092, 283.1492, 284.1492, 
    284.6392, 283.4292, 284.1592, 284.7492, 285.1892, 285.1292, 284.2492, 
    282.4292, 281.2392, 281.8892, 283.2292, 284.2292, 284.7192, 283.5092, 
    284.2392, 284.8292, 285.2692, 285.2092, 284.3292, 282.5092, 281.3192, 
    281.9692, 283.3092, 284.3092, 284.7992, 283.5492, 284.2792, 284.8692, 
    285.3092, 285.2492, 284.3692, 282.5492, 281.3592, 282.0092, 283.3492, 
    284.3492, 284.8392, 283.5892, 284.3192, 284.9092, 285.3492, 285.2892, 
    284.4092, 282.5892, 281.3992, 282.0492, 283.3892, 284.3892, 284.8792, 
    283.6292, 284.3592, 284.9492, 285.3892, 285.3292, 284.4492, 282.6292, 
    281.4392, 282.0892, 283.4292, 284.4292, 284.9192, 283.6692, 284.3992, 
    284.9892, 285.4292, 285.3692, 284.4892, 282.6692, 281.4792, 282.1292, 
    283.4692, 284.4692, 284.9592, 283.7092, 284.4392, 285.0292, 285.4692, 
    285.4092, 284.5292, 282.7092, 281.5192, 282.1692, 283.5092, 284.5092, 
    284.9992, 283.7492, 284.4792, 285.0692, 285.5092, 285.4492, 284.5692, 
    282.7492, 281.5592, 282.2092, 283.5492, 284.5492, 285.0392, 283.7892, 
    284.5192, 285.1092, 285.5492, 285.4892, 284.6092, 282.7892, 281.5992, 
    282.2492, 283.5892, 284.5892, 285.0792, 283.8292, 284.5592, 285.1492, 
    285.5892, 285.5292, 284.6492, 282.8292, 281.6392, 282.2892, 283.6292, 
    284.6292, 285.1192, 283.8692, 284.5992, 285.1892, 285.6292, 285.5692, 
    284.6892, 282.8692, 281.6792, 282.3292, 283.6692, 284.6692, 285.1592, 
    283.9092, 284.6392, 285.2292, 285.6692, 285.6092, 284.7292, 282.9092, 
    281.7192, 282.3692, 283.7092, 284.7092, 285.1992, 283.9292, 284.6592, 
    285.2492, 285.6892, 285.6292, 284.7492, 282.9292, 281.7392, 282.3892, 
    283.7292, 284.7292, 285.2192, 283.9492, 284.6792, 285.2692, 285.7092, 
    285.6492, 284.7692, 282.9492, 281.7592, 282.4092, 283.7492, 284.7492, 
    285.2392, 283.9692, 284.6992, 285.2892, 285.7292, 285.6692, 284.7892, 
    282.9692, 281.7792, 282.4292, 283.7692, 284.7692, 285.2592, 283.9892, 
    284.7192, 285.3092, 285.7492, 285.6892, 284.8092, 282.9892, 281.7992, 
    282.4492, 283.7892, 284.7892, 285.2792, 284.0092, 284.7392, 285.3292, 
    285.7692, 285.7092, 284.8292, 283.0092, 281.8192, 282.4692, 283.8092, 
    284.8092, 285.2992, 284.0292, 284.7592, 285.3492, 285.7892, 285.7292, 
    284.8492, 283.0292, 281.8392, 282.4892, 283.8292, 284.8292, 285.3192, 
    284.0492, 284.7792, 285.3692, 285.8092, 285.7492, 284.8692, 283.0492, 
    281.8592, 282.5092, 283.8492, 284.8492, 285.3392, 284.0692, 284.7992, 
    285.3892, 285.8292, 285.7692, 284.8892, 283.0692, 281.8792, 282.5292, 
    283.8692, 284.8692, 285.3592, 284.0892, 284.8192, 285.4092, 285.8492, 
    285.7892, 284.9092, 283.0892, 281.8992, 282.5492, 283.8892, 284.8892, 
    285.3792, 284.1092, 284.8392, 285.4292, 285.8692, 285.8092, 284.9292, 
    283.1092, 281.9192, 282.5692, 283.9092, 284.9092, 285.3992, 283.9892, 
    284.7192, 285.3092, 285.7492, 285.6892, 284.8092, 282.9892, 281.7992, 
    282.4492, 283.7892, 284.7892, 285.2792, 283.8692, 284.5992, 285.1892, 
    285.6292, 285.5692, 284.6892, 282.8692, 281.6792, 282.3292, 283.6692, 
    284.6692, 285.1592, 283.7492, 284.4792, 285.0692, 285.5092, 285.4492, 
    284.5692, 282.7492, 281.5592, 282.2092, 283.5492, 284.5492, 285.0392, 
    283.6292, 284.3592, 284.9492, 285.3892, 285.3292, 284.4492, 282.6292, 
    281.4392, 282.0892, 283.4292, 284.4292, 284.9192, 283.5092, 284.2392, 
    284.8292, 285.2692, 285.2092, 284.3292, 282.5092, 281.3192, 281.9692, 
    283.3092, 284.3092, 284.7992, 283.4292, 284.1592, 284.7492, 285.1892, 
    285.1292, 284.2492, 282.4292, 281.2392, 281.8892, 283.2292, 284.2292, 
    284.7192, 283.3492, 284.0792, 284.6692, 285.1092, 285.0492, 284.1692, 
    282.3492, 281.1592, 281.8092, 283.1492, 284.1492, 284.6392, 283.2692, 
    283.9992, 284.5892, 285.0292, 284.9692, 284.0892, 282.2692, 281.0792, 
    281.7292, 283.0692, 284.0692, 284.5592, 283.1892, 283.9192, 284.5092, 
    284.9492, 284.8892, 284.0092, 282.1892, 280.9992, 281.6492, 282.9892, 
    283.9892, 284.4792, 283.1092, 283.8392, 284.4292, 284.8692, 284.8092, 
    283.9292, 282.1092, 280.9192, 281.5692, 282.9092, 283.9092, 284.3992, 
    283.2092, 283.9392, 284.5292, 284.9692, 284.9092, 284.0292, 282.2092, 
    281.0192, 281.6692, 283.0092, 284.0092, 284.4992, 283.3092, 284.0392, 
    284.6292, 285.0692, 285.0092, 284.1292, 282.3092, 281.1192, 281.7692, 
    283.1092, 284.1092, 284.5992, 283.4092, 284.1392, 284.7292, 285.1692, 
    285.1092, 284.2292, 282.4092, 281.2192, 281.8692, 283.2092, 284.2092, 
    284.6992, 283.5092, 284.2392, 284.8292, 285.2692, 285.2092, 284.3292, 
    282.5092, 281.3192, 281.9692, 283.3092, 284.3092, 284.7992, 283.6092, 
    284.3392, 284.9292, 285.3692, 285.3092, 284.4292, 282.6092, 281.4192, 
    282.0692, 283.4092, 284.4092, 284.8992, 283.7692, 284.4992, 285.0892, 
    285.5292, 285.4692, 284.5892, 282.7692, 281.5792, 282.2292, 283.5692, 
    284.5692, 285.0592, 283.9292, 284.6592, 285.2492, 285.6892, 285.6292, 
    284.7492, 282.9292, 281.7392, 282.3892, 283.7292, 284.7292, 285.2192, 
    284.0892, 284.8192, 285.4092, 285.8492, 285.7892, 284.9092, 283.0892, 
    281.8992, 282.5492, 283.8892, 284.8892, 285.3792, 284.2492, 284.9792, 
    285.5692, 286.0092, 285.9492, 285.0692, 283.2492, 282.0592, 282.7092, 
    284.0492, 285.0492, 285.5392, 284.4092, 285.1392, 285.7292, 286.1692, 
    286.1092, 285.2292, 283.4092, 282.2192, 282.8692, 284.2092, 285.2092, 
    285.6992, 284.5492, 285.2792, 285.8692, 286.3092, 286.2492, 285.3692, 
    283.5492, 282.3592, 283.0092, 284.3492, 285.3492, 285.8392, 284.6892, 
    285.4192, 286.0092, 286.4492, 286.3892, 285.5092, 283.6892, 282.4992, 
    283.1492, 284.4892, 285.4892, 285.9792, 284.8292, 285.5592, 286.1492, 
    286.5892, 286.5292, 285.6492, 283.8292, 282.6392, 283.2892, 284.6292, 
    285.6292, 286.1192, 284.9692, 285.6992, 286.2892, 286.7292, 286.6692, 
    285.7892, 283.9692, 282.7792, 283.4292, 284.7692, 285.7692, 286.2592, 
    285.1092, 285.8392, 286.4292, 286.8692, 286.8092, 285.9292, 284.1092, 
    282.9192, 283.5692, 284.9092, 285.9092, 286.3992, 285.2692, 285.9992, 
    286.5892, 287.0292, 286.9692, 286.0892, 284.2692, 283.0792, 283.7292, 
    285.0692, 286.0692, 286.5592, 285.4292, 286.1592, 286.7492, 287.1892, 
    287.1292, 286.2492, 284.4292, 283.2392, 283.8892, 285.2292, 286.2292, 
    286.7192, 285.5892, 286.3192, 286.9092, 287.3492, 287.2892, 286.4092, 
    284.5892, 283.3992, 284.0492, 285.3892, 286.3892, 286.8792, 285.7492, 
    286.4792, 287.0692, 287.5092, 287.4492, 286.5692, 284.7492, 283.5592, 
    284.2092, 285.5492, 286.5492, 287.0392, 285.9092, 286.6392, 287.2292, 
    287.6692, 287.6092, 286.7292, 284.9092, 283.7192, 284.3692, 285.7092, 
    286.7092, 287.1992, 286.0492, 286.7792, 287.3692, 287.8092, 287.7492, 
    286.8692, 285.0492, 283.8592, 284.5092, 285.8492, 286.8492, 287.3392, 
    286.1892, 286.9192, 287.5092, 287.9492, 287.8892, 287.0092, 285.1892, 
    283.9992, 284.6492, 285.9892, 286.9892, 287.4792, 286.3292, 287.0592, 
    287.6492, 288.0892, 288.0292, 287.1492, 285.3292, 284.1392, 284.7892, 
    286.1292, 287.1292, 287.6192, 286.4692, 287.1992, 287.7892, 288.2292, 
    288.1692, 287.2892, 285.4692, 284.2792, 284.9292, 286.2692, 287.2692, 
    287.7592, 286.6092, 287.3392, 287.9292, 288.3692, 288.3092, 287.4292, 
    285.6092, 284.4192, 285.0692, 286.4092, 287.4092, 287.8992, 286.7292, 
    287.4592, 288.0492, 288.4892, 288.4292, 287.5492, 285.7292, 284.5392, 
    285.1892, 286.5292, 287.5292, 288.0192, 286.8492, 287.5792, 288.1692, 
    288.6092, 288.5492, 287.6692, 285.8492, 284.6592, 285.3092, 286.6492, 
    287.6492, 288.1392, 286.9692, 287.6992, 288.2892, 288.7292, 288.6692, 
    287.7892, 285.9692, 284.7792, 285.4292, 286.7692, 287.7692, 288.2592, 
    287.0892, 287.8192, 288.4092, 288.8492, 288.7892, 287.9092, 286.0892, 
    284.8992, 285.5492, 286.8892, 287.8892, 288.3792, 287.2092, 287.9392, 
    288.5292, 288.9692, 288.9092, 288.0292, 286.2092, 285.0192, 285.6692, 
    287.0092, 288.0092, 288.4992, 287.4492, 288.1792, 288.7692, 289.2092, 
    289.1492, 288.2692, 286.4492, 285.2592, 285.9092, 287.2492, 288.2492, 
    288.7392, 287.6892, 288.4192, 289.0092, 289.4492, 289.3892, 288.5092, 
    286.6892, 285.4992, 286.1492, 287.4892, 288.4892, 288.9792, 287.9292, 
    288.6592, 289.2492, 289.6892, 289.6292, 288.7492, 286.9292, 285.7392, 
    286.3892, 287.7292, 288.7292, 289.2192, 288.1692, 288.8992, 289.4892, 
    289.9292, 289.8692, 288.9892, 287.1692, 285.9792, 286.6292, 287.9692, 
    288.9692, 289.4592, 288.4092, 289.1392, 289.7292, 290.1692, 290.1092, 
    289.2292, 287.4092, 286.2192, 286.8692, 288.2092, 289.2092, 289.6992, 
    288.8092, 289.5392, 290.1292, 290.5692, 290.5092, 289.6292, 287.8092, 
    286.6192, 287.2692, 288.6092, 289.6092, 290.0992, 289.2092, 289.9392, 
    290.5292, 290.9692, 290.9092, 290.0292, 288.2092, 287.0192, 287.6692, 
    289.0092, 290.0092, 290.4992, 289.6092, 290.3392, 290.9292, 291.3692, 
    291.3092, 290.4292, 288.6092, 287.4192, 288.0692, 289.4092, 290.4092, 
    290.8992, 290.0092, 290.7392, 291.3292, 291.7692, 291.7092, 290.8292, 
    289.0092, 287.8192, 288.4692, 289.8092, 290.8092, 291.2992, 290.4092, 
    291.1392, 291.7292, 292.1692, 292.1092, 291.2292, 289.4092, 288.2192, 
    288.8692, 290.2092, 291.2092, 291.6992, 290.8692, 291.5992, 292.1892, 
    292.6292, 292.5692, 291.6892, 289.8692, 288.6792, 289.3292, 290.6692, 
    291.6692, 292.1592, 291.3292, 292.0592, 292.6492, 293.0892, 293.0292, 
    292.1492, 290.3292, 289.1392, 289.7892, 291.1292, 292.1292, 292.6192, 
    291.7892, 292.5192, 293.1092, 293.5492, 293.4892, 292.6092, 290.7892, 
    289.5992, 290.2492, 291.5892, 292.5892, 293.0792, 292.2492, 292.9792, 
    293.5692, 294.0092, 293.9492, 293.0692, 291.2492, 290.0592, 290.7092, 
    292.0492, 293.0492, 293.5392, 292.7092, 293.4392, 294.0292, 294.4692, 
    294.4092, 293.5292, 291.7092, 290.5192, 291.1692, 292.5092, 293.5092, 
    293.9992, 292.9492, 293.6792, 294.2692, 294.7092, 294.6492, 293.7692, 
    291.9492, 290.7592, 291.4092, 292.7492, 293.7492, 294.2392, 293.1892, 
    293.9192, 294.5092, 294.9492, 294.8892, 294.0092, 292.1892, 290.9992, 
    291.6492, 292.9892, 293.9892, 294.4792, 293.4292, 294.1592, 294.7492, 
    295.1892, 295.1292, 294.2492, 292.4292, 291.2392, 291.8892, 293.2292, 
    294.2292, 294.7192, 293.6692, 294.3992, 294.9892, 295.4292, 295.3692, 
    294.4892, 292.6692, 291.4792, 292.1292, 293.4692, 294.4692, 294.9592, 
    293.9092, 294.6392, 295.2292, 295.6692, 295.6092, 294.7292, 292.9092, 
    291.7192, 292.3692, 293.7092, 294.7092, 295.1992, 294.0292, 294.7592, 
    295.3492, 295.7892, 295.7292, 294.8492, 293.0292, 291.8392, 292.4892, 
    293.8292, 294.8292, 295.3192, 294.1492, 294.8792, 295.4692, 295.9092, 
    295.8492, 294.9692, 293.1492, 291.9592, 292.6092, 293.9492, 294.9492, 
    295.4392, 294.2692, 294.9992, 295.5892, 296.0292, 295.9692, 295.0892, 
    293.2692, 292.0792, 292.7292, 294.0692, 295.0692, 295.5592, 294.3892, 
    295.1192, 295.7092, 296.1492, 296.0892, 295.2092, 293.3892, 292.1992, 
    292.8492, 294.1892, 295.1892, 295.6792, 294.5092, 295.2392, 295.8292, 
    296.2692, 296.2092, 295.3292, 293.5092, 292.3192, 292.9692, 294.3092, 
    295.3092, 295.7992, 294.7092, 295.4392, 296.0292, 296.4692, 296.4092, 
    295.5292, 293.7092, 292.5192, 293.1692, 294.5092, 295.5092, 295.9992, 
    294.9092, 295.6392, 296.2292, 296.6692, 296.6092, 295.7292, 293.9092, 
    292.7192, 293.3692, 294.7092, 295.7092, 296.1992, 295.1092, 295.8392, 
    296.4292, 296.8692, 296.8092, 295.9292, 294.1092, 292.9192, 293.5692, 
    294.9092, 295.9092, 296.3992, 295.3092, 296.0392, 296.6292, 297.0692, 
    297.0092, 296.1292, 294.3092, 293.1192, 293.7692, 295.1092, 296.1092, 
    296.5992, 295.5092, 296.2392, 296.8292, 297.2692, 297.2092, 296.3292, 
    294.5092, 293.3192, 293.9692, 295.3092, 296.3092, 296.7992, 295.8692, 
    296.5992, 297.1892, 297.6292, 297.5692, 296.6892, 294.8692, 293.6792, 
    294.3292, 295.6692, 296.6692, 297.1592, 296.2292, 296.9592, 297.5492, 
    297.9892, 297.9292, 297.0492, 295.2292, 294.0392, 294.6892, 296.0292, 
    297.0292, 297.5192, 296.5892, 297.3192, 297.9092, 298.3492, 298.2892, 
    297.4092, 295.5892, 294.3992, 295.0492, 296.3892, 297.3892, 297.8792, 
    296.9492, 297.6792, 298.2692, 298.7092, 298.6492, 297.7692, 295.9492, 
    294.7592, 295.4092, 296.7492, 297.7492, 298.2392, 297.3092, 298.0392, 
    298.6292, 299.0692, 299.0092, 298.1292, 296.3092, 295.1192, 295.7692, 
    297.1092, 298.1092, 298.5992, 297.7292, 298.4592, 299.0492, 299.4892, 
    299.4292, 298.5492, 296.7292, 295.5392, 296.1892, 297.5292, 298.5292, 
    299.0192, 298.1492, 298.8792, 299.4692, 299.9092, 299.8492, 298.9692, 
    297.1492, 295.9592, 296.6092, 297.9492, 298.9492, 299.4392, 298.5692, 
    299.2992, 299.8892, 300.3292, 300.2692, 299.3892, 297.5692, 296.3792, 
    297.0292, 298.3692, 299.3692, 299.8592, 298.9892, 299.7192, 300.3092, 
    300.7492, 300.6892, 299.8092, 297.9892, 296.7992, 297.4492, 298.7892, 
    299.7892, 300.2792, 299.4092, 300.1392, 300.7292, 301.1692, 301.1092, 
    300.2292, 298.4092, 297.2192, 297.8692, 299.2092, 300.2092, 300.6992, 
    299.7492, 300.4792, 301.0692, 301.5092, 301.4492, 300.5692, 298.7492, 
    297.5592, 298.2092, 299.5492, 300.5492, 301.0392, 300.0892, 300.8192, 
    301.4092, 301.8492, 301.7892, 300.9092, 299.0892, 297.8992, 298.5492, 
    299.8892, 300.8892, 301.3792, 300.4292, 301.1592, 301.7492, 302.1892, 
    302.1292, 301.2492, 299.4292, 298.2392, 298.8892, 300.2292, 301.2292, 
    301.7192, 300.7692, 301.4992, 302.0892, 302.5292, 302.4692, 301.5892, 
    299.7692, 298.5792, 299.2292, 300.5692, 301.5692, 302.0592, 301.1092, 
    301.8392, 302.4292, 302.8692, 302.8092, 301.9292, 300.1092, 298.9192, 
    299.5692, 300.9092, 301.9092, 302.3992, 301.4292, 302.1592, 302.7492, 
    303.1892, 303.1292, 302.2492, 300.4292, 299.2392, 299.8892, 301.2292, 
    302.2292, 302.7192, 301.7492, 302.4792, 303.0692, 303.5092, 303.4492, 
    302.5692, 300.7492, 299.5592, 300.2092, 301.5492, 302.5492, 303.0392, 
    302.0692, 302.7992, 303.3892, 303.8292, 303.7692, 302.8892, 301.0692, 
    299.8792, 300.5292, 301.8692, 302.8692, 303.3592, 302.3892, 303.1192, 
    303.7092, 304.1492, 304.0892, 303.2092, 301.3892, 300.1992, 300.8492, 
    302.1892, 303.1892, 303.6792, 302.7092, 303.4392, 304.0292, 304.4692, 
    304.4092, 303.5292, 301.7092, 300.5192, 301.1692, 302.5092, 303.5092, 
    303.9992, 303.1092, 303.8392, 304.4292, 304.8692, 304.8092, 303.9292, 
    302.1092, 300.9192, 301.5692, 302.9092, 303.9092, 304.3992, 303.5092, 
    304.2392, 304.8292, 305.2692, 305.2092, 304.3292, 302.5092, 301.3192, 
    301.9692, 303.3092, 304.3092, 304.7992, 303.9092, 304.6392, 305.2292, 
    305.6692, 305.6092, 304.7292, 302.9092, 301.7192, 302.3692, 303.7092, 
    304.7092, 305.1992, 304.3092, 305.0392, 305.6292, 306.0692, 306.0092, 
    305.1292, 303.3092, 302.1192, 302.7692, 304.1092, 305.1092, 305.5992, 
    304.7092, 305.4392, 306.0292, 306.4692, 306.4092, 305.5292, 303.7092, 
    302.5192, 303.1692, 304.5092, 305.5092, 305.9992, 305.1492, 305.8792, 
    306.4692, 306.9092, 306.8492, 305.9692, 304.1492, 302.9592, 303.6092, 
    304.9492, 305.9492, 306.4392, 305.5892, 306.3192, 306.9092, 307.3492, 
    307.2892, 306.4092, 304.5892, 303.3992, 304.0492, 305.3892, 306.3892, 
    306.8792, 306.0292, 306.7592, 307.3492, 307.7892, 307.7292, 306.8492, 
    305.0292, 303.8392, 304.4892, 305.8292, 306.8292, 307.3192, 306.4692, 
    307.1992, 307.7892, 308.2292, 308.1692, 307.2892, 305.4692, 304.2792, 
    304.9292, 306.2692, 307.2692, 307.7592, 306.9092, 307.6392, 308.2292, 
    308.6692, 308.6092, 307.7292, 305.9092, 304.7192, 305.3692, 306.7092, 
    307.7092, 308.1992, 307.3492, 308.0792, 308.6692, 309.1092, 309.0492, 
    308.1692, 306.3492, 305.1592, 305.8092, 307.1492, 308.1492, 308.6392, 
    307.7892, 308.5192, 309.1092, 309.5492, 309.4892, 308.6092, 306.7892, 
    305.5992, 306.2492, 307.5892, 308.5892, 309.0792, 308.2292, 308.9592, 
    309.5492, 309.9892, 309.9292, 309.0492, 307.2292, 306.0392, 306.6892, 
    308.0292, 309.0292, 309.5192, 308.6692, 309.3992, 309.9892, 310.4292, 
    310.3692, 309.4892, 307.6692, 306.4792, 307.1292, 308.4692, 309.4692, 
    309.9592, 309.1092, 309.8392, 310.4292, 310.8692, 310.8092, 309.9292, 
    308.1092, 306.9192, 307.5692, 308.9092, 309.9092, 310.3992, 309.3092, 
    310.0392, 310.6292, 311.0692, 311.0092, 310.1292, 308.3092, 307.1192, 
    307.7692, 309.1092, 310.1092, 310.5992, 309.5092, 310.2392, 310.8292, 
    311.2692, 311.2092, 310.3292, 308.5092, 307.3192, 307.9692, 309.3092, 
    310.3092, 310.7992, 309.7092, 310.4392, 311.0292, 311.4692, 311.4092, 
    310.5292, 308.7092, 307.5192, 308.1692, 309.5092, 310.5092, 310.9992, 
    309.9092, 310.6392, 311.2292, 311.6692, 311.6092, 310.7292, 308.9092, 
    307.7192, 308.3692, 309.7092, 310.7092, 311.1992, 310.1092, 310.8392, 
    311.4292, 311.8692, 311.8092, 310.9292, 309.1092, 307.9192, 308.5692, 
    309.9092, 310.9092, 311.3992, 310.0492, 310.7792, 311.3692, 311.8092, 
    311.7492, 310.8692, 309.0492, 307.8592, 308.5092, 309.8492, 310.8492, 
    311.3392, 309.9892, 310.7192, 311.3092, 311.7492, 311.6892, 310.8092, 
    308.9892, 307.7992, 308.4492, 309.7892, 310.7892, 311.2792, 309.9292, 
    310.6592, 311.2492, 311.6892, 311.6292, 310.7492, 308.9292, 307.7392, 
    308.3892, 309.7292, 310.7292, 311.2192, 309.8692, 310.5992, 311.1892, 
    311.6292, 311.5692, 310.6892, 308.8692, 307.6792, 308.3292, 309.6692, 
    310.6692, 311.1592, 309.8092, 310.5392, 311.1292, 311.5692, 311.5092, 
    310.6292, 308.8092, 307.6192, 308.2692, 309.6092, 310.6092, 311.0992, 
    309.9292, 310.6592, 311.2492, 311.6892, 311.6292, 310.7492, 308.9292, 
    307.7392, 308.3892, 309.7292, 310.7292, 311.2192, 310.0492, 310.7792, 
    311.3692, 311.8092, 311.7492, 310.8692, 309.0492, 307.8592, 308.5092, 
    309.8492, 310.8492, 311.3392, 310.1692, 310.8992, 311.4892, 311.9292, 
    311.8692, 310.9892, 309.1692, 307.9792, 308.6292, 309.9692, 310.9692, 
    311.4592, 310.2892, 311.0192, 311.6092, 312.0492, 311.9892, 311.1092, 
    309.2892, 308.0992, 308.7492, 310.0892, 311.0892, 311.5792, 310.4092, 
    311.1392, 311.7292, 312.1692, 312.1092, 311.2292, 309.4092, 308.2192, 
    308.8692, 310.2092, 311.2092, 311.6992, 310.8692, 311.5992, 312.1892, 
    312.6292, 312.5692, 311.6892, 309.8692, 308.6792, 309.3292, 310.6692, 
    311.6692, 312.1592, 311.3292, 312.0592, 312.6492, 313.0892, 313.0292, 
    312.1492, 310.3292, 309.1392, 309.7892, 311.1292, 312.1292, 312.6192, 
    311.7892, 312.5192, 313.1092, 313.5492, 313.4892, 312.6092, 310.7892, 
    309.5992, 310.2492, 311.5892, 312.5892, 313.0792, 312.2492, 312.9792, 
    313.5692, 314.0092, 313.9492, 313.0692, 311.2492, 310.0592, 310.7092, 
    312.0492, 313.0492, 313.5392, 312.7092, 313.4392, 314.0292, 314.4692, 
    314.4092, 313.5292, 311.7092, 310.5192, 311.1692, 312.5092, 313.5092, 
    313.9992, 313.4542, 314.1842, 314.7742, 315.2142, 315.1542, 314.2742, 
    312.4542, 311.2642, 311.9142, 313.2542, 314.2542, 314.7442, 314.1992, 
    314.9292, 315.5192, 315.9592, 315.8992, 315.0192, 313.1992, 312.0092, 
    312.6592, 313.9992, 314.9992, 315.4892, 314.9442, 315.6742, 316.2642, 
    316.7042, 316.6442, 315.7642, 313.9442, 312.7542, 313.4042, 314.7442, 
    315.7442, 316.2342, 315.6892, 316.4192, 317.0092, 317.4492, 317.3892, 
    316.5092, 314.6892, 313.4992, 314.1492, 315.4892, 316.4892, 316.9792, 
    316.6192, 317.3492, 317.9392, 318.3792, 318.3192, 317.4392, 315.6192, 
    314.4292, 315.0792, 316.4192, 317.4192, 317.9092, 317.3492, 318.0792, 
    318.6692, 319.1092, 319.0492, 318.1692, 316.3492, 315.1592, 315.8092, 
    317.1492, 318.1492, 318.6392, 318.1592, 318.8892, 319.4792, 319.9192, 
    319.8592, 318.9792, 317.1592, 315.9692, 316.6192, 317.9592, 318.9592, 
    319.4492, 318.6992, 319.4292, 320.0192, 320.4592, 320.3992, 319.5192, 
    317.6992, 316.5092, 317.1592, 318.4992, 319.4992, 319.9892, 319.3292, 
    320.0592, 320.6492, 321.0892, 321.0292, 320.1492, 318.3292, 317.1392, 
    317.7892, 319.1292, 320.1292, 320.6192, 319.7492, 320.4792, 321.0692, 
    321.5092, 321.4492, 320.5692, 318.7492, 317.5592, 318.2092, 319.5492, 
    320.5492, 321.0392, 321.0792, 321.8092, 322.3992, 322.8392, 322.7792, 
    321.8992, 320.0792, 318.8892, 319.5392, 320.8792, 321.8792, 322.3692, 
    321.8892, 322.6192, 323.2092, 323.6492, 323.5892, 322.7092, 320.8892, 
    319.6992, 320.3492, 321.6892, 322.6892, 323.1792, 322.7592, 323.4892, 
    324.0792, 324.5192, 324.4592, 323.5792, 321.7592, 320.5692, 321.2192, 
    322.5592, 323.5592, 324.0492, 324.3292, 325.0592, 325.6492, 326.0892, 
    326.0292, 325.1492, 323.3292, 322.1392, 322.7892, 324.1292, 325.1292, 
    325.6192, 325.3892, 326.1192, 326.7092, 327.1492, 327.0892, 326.2092, 
    324.3892, 323.1992, 323.8492, 325.1892, 326.1892, 326.6792, 326.0292, 
    326.7592, 327.3492, 327.7892, 327.7292, 326.8492, 325.0292, 323.8392, 
    324.4892, 325.8292, 326.8292, 327.3192, 327.1692, 327.8992, 328.4892, 
    328.9292, 328.8692, 327.9892, 326.1692, 324.9792, 325.6292, 326.9692, 
    327.9692, 328.4592, 329.3892, 330.1192, 330.7092, 331.1492, 331.0892, 
    330.2092, 328.3892, 327.1992, 327.8492, 329.1892, 330.1892, 330.6792, 
    329.8992, 330.6292, 331.2192, 331.6592, 331.5992, 330.7192, 328.8992, 
    327.7092, 328.3592, 329.6992, 330.6992, 331.1892, 330.8392, 331.5692, 
    332.1592, 332.5992, 332.5392, 331.6592, 329.8392, 328.6492, 329.2992, 
    330.6392, 331.6392, 332.1292, 331.7392, 332.4692, 333.0592, 333.4992, 
    333.4392, 332.5592, 330.7392, 329.5492, 330.1992, 331.5392, 332.5392, 
    333.0292, 333.5492, 334.2792, 334.8692, 335.3092, 335.2492, 334.3692, 
    332.5492, 331.3592, 332.0092, 333.3492, 334.3492, 334.8392, 335.1192, 
    335.8492, 336.4392, 336.8792, 336.8192, 335.9392, 334.1192, 332.9292, 
    333.5792, 334.9192, 335.9192, 336.4092, 336.5492, 337.2792, 337.8692, 
    338.3092, 338.2492, 337.3692, 335.5492, 334.3592, 335.0092, 336.3492, 
    337.3492, 337.8392, 338.4, 339.11, 339.44, 339.84, 340.29, 339.84, 
    338.29, 337.06, 336.9, 337.68, 338.78, 339.49, 340.1892, 340.7592, 
    341.3892, 341.6892, 341.4392, 340.6392, 339.2292, 338.0892, 337.9892, 
    339.0792, 340.1892, 340.7592, 341.9942, 342.5742, 342.8542, 343.1442, 
    342.9842, 342.1142, 340.3742, 338.7342, 338.7842, 340.2342, 341.5742, 
    342.3942, 342.99, 343.36, 343.66, 344.13, 344.46, 344.12, 342.76, 341.24, 
    341.15, 342.37, 343.45, 344.11, 345.1167, 345.6167, 345.7567, 345.9867, 
    346.1267, 345.3667, 343.9967, 343.0067, 342.9267, 343.7867, 344.9567, 
    345.7967, 346.1625, 346.6125, 347.4525, 347.7525, 347.5925, 347.0725, 
    345.7325, 344.2225, 344.1825, 345.4525, 346.6025, 347.3625, 347.7517, 
    347.9817, 348.3517, 348.8617, 348.9617, 348.4017, 346.9317, 345.5617, 
    345.5017, 346.6717, 347.9417, 348.4017, 348.6467, 349.1967, 349.9167, 
    350.6067, 350.8867, 350.1067, 348.4867, 347.2367, 347.3267, 348.5967, 
    349.8767, 350.8367, 351.4408, 352.0008, 352.3808, 352.8308, 352.9908, 
    352.2908, 350.8108, 349.6308, 349.8008, 350.9708, 352.1408, 352.9908, 
    353.4225, 353.8725, 354.4225, 354.7925, 354.6025, 353.6825, 351.9725, 
    350.6225, 350.9725, 352.2625, 353.4525, 354.3225, 354.8633, 355.2733, 
    355.5933, 355.9033, 355.7933, 354.7133, 353.0933, 351.9733, 352.1833, 
    353.5833, 354.8433, 355.5833, 356.0667, 356.4967, 356.9867, 357.4967, 
    357.4167, 356.4767, 354.8367, 353.3567, 353.2367, 354.3067, 355.4667, 
    356.2567, 356.9883, 357.3383, 357.7083, 358.1983, 358.2683, 357.3183, 
    355.6283, 354.1183, 354.0283, 355.2583, 356.4383, 357.1883, 357.5867, 
    357.9167, 358.3367, 358.8067, 358.7567, 357.7167, 356.0967, 354.8167, 
    354.8467, 356.0767, 357.3267, 358.2367, 359.1133, 359.6333, 359.9933, 
    360.3433, 360.3733, 359.4333, 357.9033, 356.6833, 356.6533, 357.8933, 
    359.3233, 360.1733, 360.9283, 361.4083, 361.8783, 362.3483, 362.2683, 
    361.4083, 359.7883, 358.5283, 358.8483, 360.2183, 361.5683, 362.4483, 
    362.9475, 363.3075, 363.6275, 363.9475, 364.0975, 363.6875, 362.3775, 
    360.8775, 360.5075, 361.4775, 362.5875, 363.4375, 364.1175, 364.4675, 
    364.8575, 365.3375, 365.3475, 364.4375, 362.7675, 361.2475, 361.2375, 
    362.7775, 364.4475, 365.5175, 366.3325, 366.6025, 367.0725, 367.7225, 
    368.0025, 367.4125, 365.9825, 364.9325, 365.1825, 366.4825, 367.7425, 
    368.6125, 368.8558, 369.2558, 369.6558, 370.0358, 369.9558, 369.1058, 
    367.4358, 366.0758, 366.1958, 367.4958, 368.7858, 369.6258, 370.135, 
    370.395, 370.715, 371.095, 370.985, 370.055, 368.655, 367.505, 367.455, 
    368.655, 370.025, 370.845, 371.4367, 371.9267, 372.3367, 372.6467, 
    372.5467, 371.5967, 370.2067, 369.0667, 369.1067, 370.4567, 371.7967, 
    372.7167, 373.3767, 373.7767, 374.2467, 374.5967, 374.5767, 373.7067, 
    372.2767, 371.2167, 371.5367, 372.8167, 374.1467, 375.1267, 375.7792, 
    376.3092, 376.7492, 377.2292, 377.3892, 376.5492, 374.9992, 373.7692, 
    373.9292, 375.1992, 376.4992, 377.3592, 377.9575, 378.4775, 378.9075, 
    379.2275, 379.1475, 378.2575, 376.7075, 375.2375, 375.1375, 376.4775, 
    377.9475, 378.9175, 379.7292, 380.2692, 380.8692, 381.3192, 381.4192, 
    380.5992, 378.9392, 377.7292, 377.7592, 379.0692, 380.5292, 381.5292, 
    382.2717, 382.8917, 383.2817, 383.6117, 383.5717, 382.7017, 381.0117, 
    379.4317, 379.5717, 381.0217, 382.3817, 383.3317, 384.15, 384.67, 385.14, 
    385.4, 385.25, 384.38, 382.67, 381.41, 381.8, 383.22, 384.57, 385.58, 
    386.0392, 386.5492, 386.9592, 387.3392, 387.2992, 386.3892, 384.9092, 
    383.5792, 383.3492, 384.4792, 385.9892, 387.0792, 388.1725, 388.6225, 
    388.8525, 389.1325, 389.0925, 388.1025, 386.1525, 384.7725, 385.0725, 
    386.6425, 388.0825, 388.9825, 389.9633, 390.6733, 391.0233, 391.3233, 
    391.2933, 390.3533, 388.6933, 387.5733, 388.0433, 389.5933, 390.9633, 
    391.7033, 392.145, 392.575, 392.885, 393.265, 393.295, 392.355, 390.415, 
    389.095, 389.485, 391.045, 392.405, 393.235, 394.02, 394.61, 395.14, 
    395.4, 395.29, 394.25, 392.41, 391.3, 391.96, 393.57, 394.97, 395.8, 
    396.4125, 397.0425, 397.6325, 398.0825, 398.0925, 397.3025, 395.8125, 
    394.5725, 394.5525, 395.8525, 397.3025, 398.2225, 398.975, 399.435, 
    399.735, 400.095, 400.155, 399.185, 397.595, 396.485, 396.585, 397.845, 
    399.325, 400.305, 400.92, 401.48, 401.93, 402.32, 402.27, 401.42, 399.74, 
    398.43, 398.7, 400.16, 401.73, 403.02, 403.9633, 404.6033, 405.1933, 
    405.7033, 405.7533, 404.9633, 403.4433, 402.1233, 402.3033, 403.7533, 
    405.1033, 406.0133, 406.865, 407.455, 407.865, 408.145, 408.185, 407.395, 
    405.645, 404.115, 404.205, 405.705, 407.245, 408.295, 408.64, 409.34, 
    409.88, 410.18, 410.04, 409.17, 407.59, 406.22, 406.29, 407.76, 409.23, 
    410.3, 411.5083, 411.9283, 412.4783, 412.9183, 412.9283, 412.1183, 
    410.4683, 409.2283, 409.5083, 411.0283, 412.4583, 413.3483, 414.2267, 
    414.7467, 415.2367, 415.6567, 415.6067, 414.6767, 412.9667, 411.5267, 
    411.7967, 413.4567, 415.0467, 415.9367, 416.4767, 416.9467, 417.2367, 
    417.5567, 417.7567, 416.9467, 415.1967, 413.8967, 414.1267, 415.5767, 
    417.3267, 418.3567, 418.6675, 419.1275, 419.6475, 420.0675, 419.9375, 
    418.9175, 417.1675, 415.8975, 416.1175, 417.6275, 419.2575, 420.2875,
    419.4700, 420.3100, 420.9900, 423.3600, 424.0000, 423.6800, 421.8300,
    419.6800, 418.5000, 418.8200, 420.4600, 421.8600 ;

 N2O = 269.935, 269.945, 269.845, 269.755, 269.745, 269.795, 269.875, 
    269.935, 270.045, 270.225, 270.395, 270.505, 269.995, 270.005, 269.905, 
    269.815, 269.805, 269.855, 269.935, 269.995, 270.105, 270.285, 270.455, 
    270.565, 270.055, 270.065, 269.965, 269.875, 269.865, 269.915, 269.995, 
    270.055, 270.165, 270.345, 270.515, 270.625, 270.115, 270.125, 270.025, 
    269.935, 269.925, 269.975, 270.055, 270.115, 270.225, 270.405, 270.575, 
    270.685, 270.175, 270.185, 270.085, 269.995, 269.985, 270.035, 270.115, 
    270.175, 270.285, 270.465, 270.635, 270.745, 270.235, 270.245, 270.145, 
    270.055, 270.045, 270.095, 270.175, 270.235, 270.345, 270.525, 270.695, 
    270.805, 270.295, 270.305, 270.205, 270.115, 270.105, 270.155, 270.235, 
    270.295, 270.405, 270.585, 270.755, 270.865, 270.355, 270.365, 270.265, 
    270.175, 270.165, 270.215, 270.295, 270.355, 270.465, 270.645, 270.815, 
    270.925, 270.415, 270.425, 270.325, 270.235, 270.225, 270.275, 270.355, 
    270.415, 270.525, 270.705, 270.875, 270.985, 270.475, 270.485, 270.385, 
    270.295, 270.285, 270.335, 270.415, 270.475, 270.585, 270.765, 270.935, 
    271.045, 270.535, 270.545, 270.445, 270.355, 270.345, 270.395, 270.475, 
    270.535, 270.645, 270.825, 270.995, 271.105, 270.595, 270.605, 270.505, 
    270.415, 270.405, 270.455, 270.535, 270.595, 270.705, 270.885, 271.055, 
    271.165, 270.655, 270.665, 270.565, 270.475, 270.465, 270.515, 270.595, 
    270.655, 270.765, 270.945, 271.115, 271.225, 270.715, 270.725, 270.625, 
    270.535, 270.525, 270.575, 270.655, 270.715, 270.825, 271.005, 271.175, 
    271.285, 270.775, 270.785, 270.685, 270.595, 270.585, 270.635, 270.715, 
    270.775, 270.885, 271.065, 271.235, 271.345, 270.835, 270.845, 270.745, 
    270.655, 270.645, 270.695, 270.775, 270.835, 270.945, 271.125, 271.295, 
    271.405, 270.895, 270.905, 270.805, 270.715, 270.705, 270.755, 270.835, 
    270.895, 271.005, 271.185, 271.355, 271.465, 270.955, 270.965, 270.865, 
    270.775, 270.765, 270.815, 270.895, 270.955, 271.065, 271.245, 271.415, 
    271.525, 271.015, 271.025, 270.925, 270.835, 270.825, 270.875, 270.955, 
    271.015, 271.125, 271.305, 271.475, 271.585, 271.075, 271.085, 270.985, 
    270.895, 270.885, 270.935, 271.015, 271.075, 271.185, 271.365, 271.535, 
    271.645, 271.135, 271.145, 271.045, 270.955, 270.945, 270.995, 271.075, 
    271.135, 271.245, 271.425, 271.595, 271.705, 271.195, 271.205, 271.105, 
    271.015, 271.005, 271.055, 271.135, 271.195, 271.305, 271.485, 271.655, 
    271.765, 271.255, 271.265, 271.165, 271.075, 271.065, 271.115, 271.195, 
    271.255, 271.365, 271.545, 271.715, 271.825, 271.315, 271.325, 271.225, 
    271.135, 271.125, 271.175, 271.255, 271.315, 271.425, 271.605, 271.775, 
    271.885, 271.375, 271.385, 271.285, 271.195, 271.185, 271.235, 271.315, 
    271.375, 271.485, 271.665, 271.835, 271.945, 271.435, 271.445, 271.345, 
    271.255, 271.245, 271.295, 271.375, 271.435, 271.545, 271.725, 271.895, 
    272.005, 271.495, 271.505, 271.405, 271.315, 271.305, 271.355, 271.435, 
    271.495, 271.605, 271.785, 271.955, 272.065, 271.555, 271.565, 271.465, 
    271.375, 271.365, 271.415, 271.495, 271.555, 271.665, 271.845, 272.015, 
    272.125, 271.615, 271.625, 271.525, 271.435, 271.425, 271.475, 271.555, 
    271.615, 271.725, 271.905, 272.075, 272.185, 271.675, 271.685, 271.585, 
    271.495, 271.485, 271.535, 271.615, 271.675, 271.785, 271.965, 272.135, 
    272.245, 271.735, 271.745, 271.645, 271.555, 271.545, 271.595, 271.675, 
    271.735, 271.845, 272.025, 272.195, 272.305, 271.795, 271.805, 271.705, 
    271.615, 271.605, 271.655, 271.735, 271.795, 271.905, 272.085, 272.255, 
    272.365, 271.855, 271.865, 271.765, 271.675, 271.665, 271.715, 271.795, 
    271.855, 271.965, 272.145, 272.315, 272.425, 271.915, 271.925, 271.825, 
    271.735, 271.725, 271.775, 271.855, 271.915, 272.025, 272.205, 272.375, 
    272.485, 271.975, 271.985, 271.885, 271.795, 271.785, 271.835, 271.915, 
    271.975, 272.085, 272.265, 272.435, 272.545, 272.035, 272.045, 271.945, 
    271.855, 271.845, 271.895, 271.975, 272.035, 272.145, 272.325, 272.495, 
    272.605, 272.095, 272.105, 272.005, 271.915, 271.905, 271.955, 272.035, 
    272.095, 272.205, 272.385, 272.555, 272.665, 272.155, 272.165, 272.065, 
    271.975, 271.965, 272.015, 272.095, 272.155, 272.265, 272.445, 272.615, 
    272.725, 272.215, 272.225, 272.125, 272.035, 272.025, 272.075, 272.155, 
    272.215, 272.325, 272.505, 272.675, 272.785, 272.275, 272.285, 272.185, 
    272.095, 272.085, 272.135, 272.215, 272.275, 272.385, 272.565, 272.735, 
    272.845, 272.335, 272.345, 272.245, 272.155, 272.145, 272.195, 272.275, 
    272.335, 272.445, 272.625, 272.795, 272.905, 272.395, 272.405, 272.305, 
    272.215, 272.205, 272.255, 272.335, 272.395, 272.505, 272.685, 272.855, 
    272.965, 272.455, 272.465, 272.365, 272.275, 272.265, 272.315, 272.395, 
    272.455, 272.565, 272.745, 272.915, 273.025, 272.515, 272.525, 272.425, 
    272.335, 272.325, 272.375, 272.455, 272.515, 272.625, 272.805, 272.975, 
    273.085, 272.575, 272.585, 272.485, 272.395, 272.385, 272.435, 272.515, 
    272.575, 272.685, 272.865, 273.035, 273.145, 272.635, 272.645, 272.545, 
    272.455, 272.445, 272.495, 272.575, 272.635, 272.745, 272.925, 273.095, 
    273.205, 272.695, 272.705, 272.605, 272.515, 272.505, 272.555, 272.635, 
    272.695, 272.805, 272.985, 273.155, 273.265, 272.755, 272.765, 272.665, 
    272.575, 272.565, 272.615, 272.695, 272.755, 272.865, 273.045, 273.215, 
    273.325, 272.815, 272.825, 272.725, 272.635, 272.625, 272.675, 272.755, 
    272.815, 272.925, 273.105, 273.275, 273.385, 272.875, 272.885, 272.785, 
    272.695, 272.685, 272.735, 272.815, 272.875, 272.985, 273.165, 273.335, 
    273.445, 272.935, 272.945, 272.845, 272.755, 272.745, 272.795, 272.875, 
    272.935, 273.045, 273.225, 273.395, 273.505, 272.983, 272.993, 272.893, 
    272.803, 272.793, 272.843, 272.923, 272.983, 273.093, 273.273, 273.443, 
    273.553, 273.031, 273.041, 272.941, 272.851, 272.841, 272.891, 272.971, 
    273.031, 273.141, 273.321, 273.491, 273.601, 273.079, 273.089, 272.989, 
    272.899, 272.889, 272.939, 273.019, 273.079, 273.189, 273.369, 273.539, 
    273.649, 273.127, 273.137, 273.037, 272.947, 272.937, 272.987, 273.067, 
    273.127, 273.237, 273.417, 273.587, 273.697, 273.175, 273.185, 273.085, 
    272.995, 272.985, 273.035, 273.115, 273.175, 273.285, 273.465, 273.635, 
    273.745, 273.223, 273.233, 273.133, 273.043, 273.033, 273.083, 273.163, 
    273.223, 273.333, 273.513, 273.683, 273.793, 273.271, 273.281, 273.181, 
    273.091, 273.081, 273.131, 273.211, 273.271, 273.381, 273.561, 273.731, 
    273.841, 273.319, 273.329, 273.229, 273.139, 273.129, 273.179, 273.259, 
    273.319, 273.429, 273.609, 273.779, 273.889, 273.367, 273.377, 273.277, 
    273.187, 273.177, 273.227, 273.307, 273.367, 273.477, 273.657, 273.827, 
    273.937, 273.415, 273.425, 273.325, 273.235, 273.225, 273.275, 273.355, 
    273.415, 273.525, 273.705, 273.875, 273.985, 273.463, 273.473, 273.373, 
    273.283, 273.273, 273.323, 273.403, 273.463, 273.573, 273.753, 273.923, 
    274.033, 273.511, 273.521, 273.421, 273.331, 273.321, 273.371, 273.451, 
    273.511, 273.621, 273.801, 273.971, 274.081, 273.559, 273.569, 273.469, 
    273.379, 273.369, 273.419, 273.499, 273.559, 273.669, 273.849, 274.019, 
    274.129, 273.607, 273.617, 273.517, 273.427, 273.417, 273.467, 273.547, 
    273.607, 273.717, 273.897, 274.067, 274.177, 273.655, 273.665, 273.565, 
    273.475, 273.465, 273.515, 273.595, 273.655, 273.765, 273.945, 274.115, 
    274.225, 273.703, 273.713, 273.613, 273.523, 273.513, 273.563, 273.643, 
    273.703, 273.813, 273.993, 274.163, 274.273, 273.751, 273.761, 273.661, 
    273.571, 273.561, 273.611, 273.691, 273.751, 273.861, 274.041, 274.211, 
    274.321, 273.799, 273.809, 273.709, 273.619, 273.609, 273.659, 273.739, 
    273.799, 273.909, 274.089, 274.259, 274.369, 273.847, 273.857, 273.757, 
    273.667, 273.657, 273.707, 273.787, 273.847, 273.957, 274.137, 274.307, 
    274.417, 273.895, 273.905, 273.805, 273.715, 273.705, 273.755, 273.835, 
    273.895, 274.005, 274.185, 274.355, 274.465, 273.943, 273.953, 273.853, 
    273.763, 273.753, 273.803, 273.883, 273.943, 274.053, 274.233, 274.403, 
    274.513, 273.991, 274.001, 273.901, 273.811, 273.801, 273.851, 273.931, 
    273.991, 274.101, 274.281, 274.451, 274.561, 274.039, 274.049, 273.949, 
    273.859, 273.849, 273.899, 273.979, 274.039, 274.149, 274.329, 274.499, 
    274.609, 274.087, 274.097, 273.997, 273.907, 273.897, 273.947, 274.027, 
    274.087, 274.197, 274.377, 274.547, 274.657, 274.135, 274.145, 274.045, 
    273.955, 273.945, 273.995, 274.075, 274.135, 274.245, 274.425, 274.595, 
    274.705, 274.183, 274.193, 274.093, 274.003, 273.993, 274.043, 274.123, 
    274.183, 274.293, 274.473, 274.643, 274.753, 274.231, 274.241, 274.141, 
    274.051, 274.041, 274.091, 274.171, 274.231, 274.341, 274.521, 274.691, 
    274.801, 274.279, 274.289, 274.189, 274.099, 274.089, 274.139, 274.219, 
    274.279, 274.389, 274.569, 274.739, 274.849, 274.327, 274.337, 274.237, 
    274.147, 274.137, 274.187, 274.267, 274.327, 274.437, 274.617, 274.787, 
    274.897, 274.375, 274.385, 274.285, 274.195, 274.185, 274.235, 274.315, 
    274.375, 274.485, 274.665, 274.835, 274.945, 274.423, 274.433, 274.333, 
    274.243, 274.233, 274.283, 274.363, 274.423, 274.533, 274.713, 274.883, 
    274.993, 274.471, 274.481, 274.381, 274.291, 274.281, 274.331, 274.411, 
    274.471, 274.581, 274.761, 274.931, 275.041, 274.519, 274.529, 274.429, 
    274.339, 274.329, 274.379, 274.459, 274.519, 274.629, 274.809, 274.979, 
    275.089, 274.567, 274.577, 274.477, 274.387, 274.377, 274.427, 274.507, 
    274.567, 274.677, 274.857, 275.027, 275.137, 274.615, 274.625, 274.525, 
    274.435, 274.425, 274.475, 274.555, 274.615, 274.725, 274.905, 275.075, 
    275.185, 274.663, 274.673, 274.573, 274.483, 274.473, 274.523, 274.603, 
    274.663, 274.773, 274.953, 275.123, 275.233, 274.711, 274.721, 274.621, 
    274.531, 274.521, 274.571, 274.651, 274.711, 274.821, 275.001, 275.171, 
    275.281, 274.759, 274.769, 274.669, 274.579, 274.569, 274.619, 274.699, 
    274.759, 274.869, 275.049, 275.219, 275.329, 274.807, 274.817, 274.717, 
    274.627, 274.617, 274.667, 274.747, 274.807, 274.917, 275.097, 275.267, 
    275.377, 274.855, 274.865, 274.765, 274.675, 274.665, 274.715, 274.795, 
    274.855, 274.965, 275.145, 275.315, 275.425, 274.903, 274.913, 274.813, 
    274.723, 274.713, 274.763, 274.843, 274.903, 275.013, 275.193, 275.363, 
    275.473, 274.951, 274.961, 274.861, 274.771, 274.761, 274.811, 274.891, 
    274.951, 275.061, 275.241, 275.411, 275.521, 274.999, 275.009, 274.909, 
    274.819, 274.809, 274.859, 274.939, 274.999, 275.109, 275.289, 275.459, 
    275.569, 275.047, 275.057, 274.957, 274.867, 274.857, 274.907, 274.987, 
    275.047, 275.157, 275.337, 275.507, 275.617, 275.095, 275.105, 275.005, 
    274.915, 274.905, 274.955, 275.035, 275.095, 275.205, 275.385, 275.555, 
    275.665, 275.143, 275.153, 275.053, 274.963, 274.953, 275.003, 275.083, 
    275.143, 275.253, 275.433, 275.603, 275.713, 275.191, 275.201, 275.101, 
    275.011, 275.001, 275.051, 275.131, 275.191, 275.301, 275.481, 275.651, 
    275.761, 275.239, 275.249, 275.149, 275.059, 275.049, 275.099, 275.179, 
    275.239, 275.349, 275.529, 275.699, 275.809, 275.287, 275.297, 275.197, 
    275.107, 275.097, 275.147, 275.227, 275.287, 275.397, 275.577, 275.747, 
    275.857, 275.335, 275.345, 275.245, 275.155, 275.145, 275.195, 275.275, 
    275.335, 275.445, 275.625, 275.795, 275.905, 275.435, 275.445, 275.345, 
    275.255, 275.245, 275.295, 275.375, 275.435, 275.545, 275.725, 275.895, 
    276.005, 275.535, 275.545, 275.445, 275.355, 275.345, 275.395, 275.475, 
    275.535, 275.645, 275.825, 275.995, 276.105, 275.635, 275.645, 275.545, 
    275.455, 275.445, 275.495, 275.575, 275.635, 275.745, 275.925, 276.095, 
    276.205, 275.735, 275.745, 275.645, 275.555, 275.545, 275.595, 275.675, 
    275.735, 275.845, 276.025, 276.195, 276.305, 275.835, 275.845, 275.745, 
    275.655, 275.645, 275.695, 275.775, 275.835, 275.945, 276.125, 276.295, 
    276.405, 275.935, 275.945, 275.845, 275.755, 275.745, 275.795, 275.875, 
    275.935, 276.045, 276.225, 276.395, 276.505, 276.035, 276.045, 275.945, 
    275.855, 275.845, 275.895, 275.975, 276.035, 276.145, 276.325, 276.495, 
    276.605, 276.135, 276.145, 276.045, 275.955, 275.945, 275.995, 276.075, 
    276.135, 276.245, 276.425, 276.595, 276.705, 276.235, 276.245, 276.145, 
    276.055, 276.045, 276.095, 276.175, 276.235, 276.345, 276.525, 276.695, 
    276.805, 276.335, 276.345, 276.245, 276.155, 276.145, 276.195, 276.275, 
    276.335, 276.445, 276.625, 276.795, 276.905, 276.435, 276.445, 276.345, 
    276.255, 276.245, 276.295, 276.375, 276.435, 276.545, 276.725, 276.895, 
    277.005, 276.535, 276.545, 276.445, 276.355, 276.345, 276.395, 276.475, 
    276.535, 276.645, 276.825, 276.995, 277.105, 276.635, 276.645, 276.545, 
    276.455, 276.445, 276.495, 276.575, 276.635, 276.745, 276.925, 277.095, 
    277.205, 276.735, 276.745, 276.645, 276.555, 276.545, 276.595, 276.675, 
    276.735, 276.845, 277.025, 277.195, 277.305, 276.835, 276.845, 276.745, 
    276.655, 276.645, 276.695, 276.775, 276.835, 276.945, 277.125, 277.295, 
    277.405, 276.935, 276.945, 276.845, 276.755, 276.745, 276.795, 276.875, 
    276.935, 277.045, 277.225, 277.395, 277.505, 277.035, 277.045, 276.945, 
    276.855, 276.845, 276.895, 276.975, 277.035, 277.145, 277.325, 277.495, 
    277.605, 277.135, 277.145, 277.045, 276.955, 276.945, 276.995, 277.075, 
    277.135, 277.245, 277.425, 277.595, 277.705, 277.235, 277.245, 277.145, 
    277.055, 277.045, 277.095, 277.175, 277.235, 277.345, 277.525, 277.695, 
    277.805, 277.335, 277.345, 277.245, 277.155, 277.145, 277.195, 277.275, 
    277.335, 277.445, 277.625, 277.795, 277.905, 277.415, 277.425, 277.325, 
    277.235, 277.225, 277.275, 277.355, 277.415, 277.525, 277.705, 277.875, 
    277.985, 277.495, 277.505, 277.405, 277.315, 277.305, 277.355, 277.435, 
    277.495, 277.605, 277.785, 277.955, 278.065, 277.575, 277.585, 277.485, 
    277.395, 277.385, 277.435, 277.515, 277.575, 277.685, 277.865, 278.035, 
    278.145, 277.655, 277.665, 277.565, 277.475, 277.465, 277.515, 277.595, 
    277.655, 277.765, 277.945, 278.115, 278.225, 277.735, 277.745, 277.645, 
    277.555, 277.545, 277.595, 277.675, 277.735, 277.845, 278.025, 278.195, 
    278.305, 277.815, 277.825, 277.725, 277.635, 277.625, 277.675, 277.755, 
    277.815, 277.925, 278.105, 278.275, 278.385, 277.895, 277.905, 277.805, 
    277.715, 277.705, 277.755, 277.835, 277.895, 278.005, 278.185, 278.355, 
    278.465, 277.975, 277.985, 277.885, 277.795, 277.785, 277.835, 277.915, 
    277.975, 278.085, 278.265, 278.435, 278.545, 278.055, 278.065, 277.965, 
    277.875, 277.865, 277.915, 277.995, 278.055, 278.165, 278.345, 278.515, 
    278.625, 278.135, 278.145, 278.045, 277.955, 277.945, 277.995, 278.075, 
    278.135, 278.245, 278.425, 278.595, 278.705, 278.235, 278.245, 278.145, 
    278.055, 278.045, 278.095, 278.175, 278.235, 278.345, 278.525, 278.695, 
    278.805, 278.335, 278.345, 278.245, 278.155, 278.145, 278.195, 278.275, 
    278.335, 278.445, 278.625, 278.795, 278.905, 278.435, 278.445, 278.345, 
    278.255, 278.245, 278.295, 278.375, 278.435, 278.545, 278.725, 278.895, 
    279.005, 278.535, 278.545, 278.445, 278.355, 278.345, 278.395, 278.475, 
    278.535, 278.645, 278.825, 278.995, 279.105, 278.635, 278.645, 278.545, 
    278.455, 278.445, 278.495, 278.575, 278.635, 278.745, 278.925, 279.095, 
    279.205, 278.715, 278.725, 278.625, 278.535, 278.525, 278.575, 278.655, 
    278.715, 278.825, 279.005, 279.175, 279.285, 278.795, 278.805, 278.705, 
    278.615, 278.605, 278.655, 278.735, 278.795, 278.905, 279.085, 279.255, 
    279.365, 278.875, 278.885, 278.785, 278.695, 278.685, 278.735, 278.815, 
    278.875, 278.985, 279.165, 279.335, 279.445, 278.955, 278.965, 278.865, 
    278.775, 278.765, 278.815, 278.895, 278.955, 279.065, 279.245, 279.415, 
    279.525, 279.035, 279.045, 278.945, 278.855, 278.845, 278.895, 278.975, 
    279.035, 279.145, 279.325, 279.495, 279.605, 279.115, 279.125, 279.025, 
    278.935, 278.925, 278.975, 279.055, 279.115, 279.225, 279.405, 279.575, 
    279.685, 279.195, 279.205, 279.105, 279.015, 279.005, 279.055, 279.135, 
    279.195, 279.305, 279.485, 279.655, 279.765, 279.275, 279.285, 279.185, 
    279.095, 279.085, 279.135, 279.215, 279.275, 279.385, 279.565, 279.735, 
    279.845, 279.355, 279.365, 279.265, 279.175, 279.165, 279.215, 279.295, 
    279.355, 279.465, 279.645, 279.815, 279.925, 279.435, 279.445, 279.345, 
    279.255, 279.245, 279.295, 279.375, 279.435, 279.545, 279.725, 279.895, 
    280.005, 279.495, 279.505, 279.405, 279.315, 279.305, 279.355, 279.435, 
    279.495, 279.605, 279.785, 279.955, 280.065, 279.555, 279.565, 279.465, 
    279.375, 279.365, 279.415, 279.495, 279.555, 279.665, 279.845, 280.015, 
    280.125, 279.615, 279.625, 279.525, 279.435, 279.425, 279.475, 279.555, 
    279.615, 279.725, 279.905, 280.075, 280.185, 279.675, 279.685, 279.585, 
    279.495, 279.485, 279.535, 279.615, 279.675, 279.785, 279.965, 280.135, 
    280.245, 279.735, 279.745, 279.645, 279.555, 279.545, 279.595, 279.675, 
    279.735, 279.845, 280.025, 280.195, 280.305, 279.835, 279.845, 279.745, 
    279.655, 279.645, 279.695, 279.775, 279.835, 279.945, 280.125, 280.295, 
    280.405, 279.935, 279.945, 279.845, 279.755, 279.745, 279.795, 279.875, 
    279.935, 280.045, 280.225, 280.395, 280.505, 280.035, 280.045, 279.945, 
    279.855, 279.845, 279.895, 279.975, 280.035, 280.145, 280.325, 280.495, 
    280.605, 280.135, 280.145, 280.045, 279.955, 279.945, 279.995, 280.075, 
    280.135, 280.245, 280.425, 280.595, 280.705, 280.235, 280.245, 280.145, 
    280.055, 280.045, 280.095, 280.175, 280.235, 280.345, 280.525, 280.695, 
    280.805, 280.375, 280.385, 280.285, 280.195, 280.185, 280.235, 280.315, 
    280.375, 280.485, 280.665, 280.835, 280.945, 280.515, 280.525, 280.425, 
    280.335, 280.325, 280.375, 280.455, 280.515, 280.625, 280.805, 280.975, 
    281.085, 280.655, 280.665, 280.565, 280.475, 280.465, 280.515, 280.595, 
    280.655, 280.765, 280.945, 281.115, 281.225, 280.795, 280.805, 280.705, 
    280.615, 280.605, 280.655, 280.735, 280.795, 280.905, 281.085, 281.255, 
    281.365, 280.935, 280.945, 280.845, 280.755, 280.745, 280.795, 280.875, 
    280.935, 281.045, 281.225, 281.395, 281.505, 281.095, 281.105, 281.005, 
    280.915, 280.905, 280.955, 281.035, 281.095, 281.205, 281.385, 281.555, 
    281.665, 281.255, 281.265, 281.165, 281.075, 281.065, 281.115, 281.195, 
    281.255, 281.365, 281.545, 281.715, 281.825, 281.415, 281.425, 281.325, 
    281.235, 281.225, 281.275, 281.355, 281.415, 281.525, 281.705, 281.875, 
    281.985, 281.575, 281.585, 281.485, 281.395, 281.385, 281.435, 281.515, 
    281.575, 281.685, 281.865, 282.035, 282.145, 281.735, 281.745, 281.645, 
    281.555, 281.545, 281.595, 281.675, 281.735, 281.845, 282.025, 282.195, 
    282.305, 281.955, 281.965, 281.865, 281.775, 281.765, 281.815, 281.895, 
    281.955, 282.065, 282.245, 282.415, 282.525, 282.175, 282.185, 282.085, 
    281.995, 281.985, 282.035, 282.115, 282.175, 282.285, 282.465, 282.635, 
    282.745, 282.395, 282.405, 282.305, 282.215, 282.205, 282.255, 282.335, 
    282.395, 282.505, 282.685, 282.855, 282.965, 282.615, 282.625, 282.525, 
    282.435, 282.425, 282.475, 282.555, 282.615, 282.725, 282.905, 283.075, 
    283.185, 282.835, 282.845, 282.745, 282.655, 282.645, 282.695, 282.775, 
    282.835, 282.945, 283.125, 283.295, 283.405, 283.055, 283.065, 282.965, 
    282.875, 282.865, 282.915, 282.995, 283.055, 283.165, 283.345, 283.515, 
    283.625, 283.275, 283.285, 283.185, 283.095, 283.085, 283.135, 283.215, 
    283.275, 283.385, 283.565, 283.735, 283.845, 283.495, 283.505, 283.405, 
    283.315, 283.305, 283.355, 283.435, 283.495, 283.605, 283.785, 283.955, 
    284.065, 283.715, 283.725, 283.625, 283.535, 283.525, 283.575, 283.655, 
    283.715, 283.825, 284.005, 284.175, 284.285, 283.935, 283.945, 283.845, 
    283.755, 283.745, 283.795, 283.875, 283.935, 284.045, 284.225, 284.395, 
    284.505, 284.135, 284.145, 284.045, 283.955, 283.945, 283.995, 284.075, 
    284.135, 284.245, 284.425, 284.595, 284.705, 284.335, 284.345, 284.245, 
    284.155, 284.145, 284.195, 284.275, 284.335, 284.445, 284.625, 284.795, 
    284.905, 284.535, 284.545, 284.445, 284.355, 284.345, 284.395, 284.475, 
    284.535, 284.645, 284.825, 284.995, 285.105, 284.735, 284.745, 284.645, 
    284.555, 284.545, 284.595, 284.675, 284.735, 284.845, 285.025, 285.195, 
    285.305, 284.935, 284.945, 284.845, 284.755, 284.745, 284.795, 284.875, 
    284.935, 285.045, 285.225, 285.395, 285.505, 285.115, 285.125, 285.025, 
    284.935, 284.925, 284.975, 285.055, 285.115, 285.225, 285.405, 285.575, 
    285.685, 285.295, 285.305, 285.205, 285.115, 285.105, 285.155, 285.235, 
    285.295, 285.405, 285.585, 285.755, 285.865, 285.475, 285.485, 285.385, 
    285.295, 285.285, 285.335, 285.415, 285.475, 285.585, 285.765, 285.935, 
    286.045, 285.655, 285.665, 285.565, 285.475, 285.465, 285.515, 285.595, 
    285.655, 285.765, 285.945, 286.115, 286.225, 285.835, 285.845, 285.745, 
    285.655, 285.645, 285.695, 285.775, 285.835, 285.945, 286.125, 286.295, 
    286.405, 285.995, 286.005, 285.905, 285.815, 285.805, 285.855, 285.935, 
    285.995, 286.105, 286.285, 286.455, 286.565, 286.155, 286.165, 286.065, 
    285.975, 285.965, 286.015, 286.095, 286.155, 286.265, 286.445, 286.615, 
    286.725, 286.315, 286.325, 286.225, 286.135, 286.125, 286.175, 286.255, 
    286.315, 286.425, 286.605, 286.775, 286.885, 286.475, 286.485, 286.385, 
    286.295, 286.285, 286.335, 286.415, 286.475, 286.585, 286.765, 286.935, 
    287.045, 286.635, 286.645, 286.545, 286.455, 286.445, 286.495, 286.575, 
    286.635, 286.745, 286.925, 287.095, 287.205, 286.855, 286.865, 286.765, 
    286.675, 286.665, 286.715, 286.795, 286.855, 286.965, 287.145, 287.315, 
    287.425, 287.075, 287.085, 286.985, 286.895, 286.885, 286.935, 287.015, 
    287.075, 287.185, 287.365, 287.535, 287.645, 287.295, 287.305, 287.205, 
    287.115, 287.105, 287.155, 287.235, 287.295, 287.405, 287.585, 287.755, 
    287.865, 287.515, 287.525, 287.425, 287.335, 287.325, 287.375, 287.455, 
    287.515, 287.625, 287.805, 287.975, 288.085, 287.735, 287.745, 287.645, 
    287.555, 287.545, 287.595, 287.675, 287.735, 287.845, 288.025, 288.195, 
    288.305, 287.975, 287.985, 287.885, 287.795, 287.785, 287.835, 287.915, 
    287.975, 288.085, 288.265, 288.435, 288.545, 288.215, 288.225, 288.125, 
    288.035, 288.025, 288.075, 288.155, 288.215, 288.325, 288.505, 288.675, 
    288.785, 288.455, 288.465, 288.365, 288.275, 288.265, 288.315, 288.395, 
    288.455, 288.565, 288.745, 288.915, 289.025, 288.695, 288.705, 288.605, 
    288.515, 288.505, 288.555, 288.635, 288.695, 288.805, 288.985, 289.155, 
    289.265, 288.935, 288.945, 288.845, 288.755, 288.745, 288.795, 288.875, 
    288.935, 289.045, 289.225, 289.395, 289.505, 289.155, 289.165, 289.065, 
    288.975, 288.965, 289.015, 289.095, 289.155, 289.265, 289.445, 289.615, 
    289.725, 289.375, 289.385, 289.285, 289.195, 289.185, 289.235, 289.315, 
    289.375, 289.485, 289.665, 289.835, 289.945, 289.595, 289.605, 289.505, 
    289.415, 289.405, 289.455, 289.535, 289.595, 289.705, 289.885, 290.055, 
    290.165, 289.815, 289.825, 289.725, 289.635, 289.625, 289.675, 289.755, 
    289.815, 289.925, 290.105, 290.275, 290.385, 290.035, 290.045, 289.945, 
    289.855, 289.845, 289.895, 289.975, 290.035, 290.145, 290.325, 290.495, 
    290.605, 290.295, 290.305, 290.205, 290.115, 290.105, 290.155, 290.235, 
    290.295, 290.405, 290.585, 290.755, 290.865, 290.555, 290.565, 290.465, 
    290.375, 290.365, 290.415, 290.495, 290.555, 290.665, 290.845, 291.015, 
    291.125, 290.815, 290.825, 290.725, 290.635, 290.625, 290.675, 290.755, 
    290.815, 290.925, 291.105, 291.275, 291.385, 291.075, 291.085, 290.985, 
    290.895, 290.885, 290.935, 291.015, 291.075, 291.185, 291.365, 291.535, 
    291.645, 291.335, 291.345, 291.245, 291.155, 291.145, 291.195, 291.275, 
    291.335, 291.445, 291.625, 291.795, 291.905, 291.635, 291.645, 291.545, 
    291.455, 291.445, 291.495, 291.575, 291.635, 291.745, 291.925, 292.095, 
    292.205, 291.935, 291.945, 291.845, 291.755, 291.745, 291.795, 291.875, 
    291.935, 292.045, 292.225, 292.395, 292.505, 292.235, 292.245, 292.145, 
    292.055, 292.045, 292.095, 292.175, 292.235, 292.345, 292.525, 292.695, 
    292.805, 292.535, 292.545, 292.445, 292.355, 292.345, 292.395, 292.475, 
    292.535, 292.645, 292.825, 292.995, 293.105, 292.835, 292.845, 292.745, 
    292.655, 292.645, 292.695, 292.775, 292.835, 292.945, 293.125, 293.295, 
    293.405, 293.235, 293.245, 293.145, 293.055, 293.045, 293.095, 293.175, 
    293.235, 293.345, 293.525, 293.695, 293.805, 293.635, 293.645, 293.545, 
    293.455, 293.445, 293.495, 293.575, 293.635, 293.745, 293.925, 294.095, 
    294.205, 294.035, 294.045, 293.945, 293.855, 293.845, 293.895, 293.975, 
    294.035, 294.145, 294.325, 294.495, 294.605, 294.435, 294.445, 294.345, 
    294.255, 294.245, 294.295, 294.375, 294.435, 294.545, 294.725, 294.895, 
    295.005, 294.835, 294.845, 294.745, 294.655, 294.645, 294.695, 294.775, 
    294.835, 294.945, 295.125, 295.295, 295.405, 295.335, 295.345, 295.245, 
    295.155, 295.145, 295.195, 295.275, 295.335, 295.445, 295.625, 295.795, 
    295.905, 295.835, 295.845, 295.745, 295.655, 295.645, 295.695, 295.775, 
    295.835, 295.945, 296.125, 296.295, 296.405, 296.335, 296.345, 296.245, 
    296.155, 296.145, 296.195, 296.275, 296.335, 296.445, 296.625, 296.795, 
    296.905, 296.835, 296.845, 296.745, 296.655, 296.645, 296.695, 296.775, 
    296.835, 296.945, 297.125, 297.295, 297.405, 297.335, 297.345, 297.245, 
    297.155, 297.145, 297.195, 297.275, 297.335, 297.445, 297.625, 297.795, 
    297.905, 297.8083, 297.8183, 297.7183, 297.6283, 297.6183, 297.6683, 
    297.7483, 297.8083, 297.9183, 298.0983, 298.2683, 298.3783, 298.2817, 
    298.2917, 298.1917, 298.1017, 298.0917, 298.1417, 298.2217, 298.2817, 
    298.3917, 298.5717, 298.7417, 298.8517, 298.755, 298.765, 298.665, 
    298.575, 298.565, 298.615, 298.695, 298.755, 298.865, 299.045, 299.215, 
    299.325, 299.975, 299.985, 299.885, 299.795, 299.785, 299.835, 299.915, 
    299.975, 300.085, 300.265, 300.435, 300.545, 300.585, 300.595, 300.495, 
    300.405, 300.395, 300.445, 300.525, 300.585, 300.695, 300.875, 301.045, 
    301.155, 301.165, 301.175, 301.075, 300.985, 300.975, 301.025, 301.105, 
    301.165, 301.275, 301.455, 301.625, 301.735, 303.495, 303.505, 303.405, 
    303.315, 303.305, 303.355, 303.435, 303.495, 303.605, 303.785, 303.955, 
    304.065, 303.715, 303.725, 303.625, 303.535, 303.525, 303.575, 303.655, 
    303.715, 303.825, 304.005, 304.175, 304.285, 303.955, 303.965, 303.865, 
    303.775, 303.765, 303.815, 303.895, 303.955, 304.065, 304.245, 304.415, 
    304.525, 304.475, 304.485, 304.385, 304.295, 304.285, 304.335, 304.415, 
    304.475, 304.585, 304.765, 304.935, 305.045, 305.305, 305.315, 305.215, 
    305.125, 305.115, 305.165, 305.245, 305.305, 305.415, 305.595, 305.765, 
    305.875, 305.485, 305.495, 305.395, 305.305, 305.295, 305.345, 305.425, 
    305.485, 305.595, 305.775, 305.945, 306.055, 306.425, 306.435, 306.335, 
    306.245, 306.235, 306.285, 306.365, 306.425, 306.535, 306.715, 306.885, 
    306.995, 307.415, 307.425, 307.325, 307.235, 307.225, 307.275, 307.355, 
    307.415, 307.525, 307.705, 307.875, 307.985, 308.715, 308.725, 308.625, 
    308.535, 308.525, 308.575, 308.655, 308.715, 308.825, 309.005, 309.175, 
    309.285, 309.505, 309.515, 309.415, 309.325, 309.315, 309.365, 309.445, 
    309.505, 309.615, 309.795, 309.965, 310.075, 309.935, 309.945, 309.845, 
    309.755, 309.745, 309.795, 309.875, 309.935, 310.045, 310.225, 310.395, 
    310.505, 310.185, 310.195, 310.095, 310.005, 309.995, 310.045, 310.125, 
    310.185, 310.295, 310.475, 310.645, 310.755, 310.915, 310.925, 310.825, 
    310.735, 310.725, 310.775, 310.855, 310.915, 311.025, 311.205, 311.375, 
    311.485, 311.715, 311.725, 311.625, 311.535, 311.525, 311.575, 311.655, 
    311.715, 311.825, 312.005, 312.175, 312.285, 312.745, 312.755, 312.655, 
    312.565, 312.555, 312.605, 312.685, 312.745, 312.855, 313.035, 313.205, 
    313.315, 313.465, 313.475, 313.375, 313.285, 313.275, 313.325, 313.405, 
    313.465, 313.575, 313.755, 313.925, 314.035, 314.135, 314.145, 314.045, 
    313.955, 313.945, 313.995, 314.075, 314.135, 314.245, 314.425, 314.595, 
    314.705, 315.085, 315.095, 314.995, 314.905, 314.895, 314.945, 315.025, 
    315.085, 315.195, 315.375, 315.545, 315.655, 316.075, 316.085, 315.985, 
    315.895, 315.885, 315.935, 316.015, 316.075, 316.185, 316.365, 316.535, 
    316.645, 316.295, 316.305, 316.205, 316.115, 316.105, 316.155, 316.235, 
    316.295, 316.405, 316.585, 316.755, 316.865, 316.9275, 316.9675, 
    316.9575, 316.8975, 316.8475, 316.8275, 316.8175, 316.8175, 316.8675, 
    316.9875, 317.1275, 317.2375, 317.2958, 317.3358, 317.4058, 317.4658, 
    317.5058, 317.5258, 317.5658, 317.6258, 317.7658, 317.9258, 318.0358, 
    318.1058, 318.175, 318.195, 318.165, 318.135, 318.135, 318.125, 318.135, 
    318.165, 318.225, 318.345, 318.555, 318.765, 318.86, 318.88, 318.86, 
    318.77, 318.65, 318.59, 318.65, 318.76, 318.89, 319.09, 319.35, 319.57, 
    319.7242, 319.8042, 319.7642, 319.6942, 319.6742, 319.6542, 319.6242, 
    319.6742, 319.8142, 319.9942, 320.1542, 320.2642, 320.3517, 320.3717, 
    320.2717, 320.1817, 320.2117, 320.2417, 320.1717, 320.2117, 320.4517, 
    320.7317, 320.9417, 321.1417, 321.3208, 321.3808, 321.3808, 321.3808, 
    321.4208, 321.4408, 321.4108, 321.3908, 321.4808, 321.6408, 321.7908, 
    321.9608, 322.2067, 322.3267, 322.2467, 322.0867, 321.9667, 321.9367, 
    322.0067, 322.1367, 322.2967, 322.4967, 322.6967, 322.8367, 322.9033, 
    322.9233, 322.9333, 322.9633, 323.0033, 323.0033, 323.0133, 323.0933, 
    323.2533, 323.5033, 323.7533, 323.9333, 324.0333, 324.0733, 324.0633, 
    324.0533, 324.0433, 324.0433, 324.0433, 324.0933, 324.2333, 324.4433, 
    324.6233, 324.7733, 324.8908, 324.9608, 324.9408, 324.9108, 324.8908, 
    324.8508, 324.8608, 324.9608, 325.1108, 325.2708, 325.4308, 325.5208, 
    325.57, 325.61, 325.67, 325.73, 325.8, 325.88, 325.94, 325.97, 326.04, 
    326.19, 326.37, 326.51, 326.6033, 326.6533, 326.7133, 326.7833, 326.8133, 
    326.8833, 327.0233, 327.1833, 327.3333, 327.5133, 327.7133, 327.8633, 
    327.9817, 328.0417, 328.0317, 327.9617, 327.9117, 327.9517, 328.0317, 
    328.1117, 328.2317, 328.4117, 328.6117, 328.7617, 328.865, 328.895, 
    328.875, 328.875, 328.895, 328.905, 328.835, 328.775, 328.855, 329.045, 
    329.225, 329.355, 329.4533, 329.5133, 329.5333, 329.5233, 329.5133, 
    329.5733, 329.6933, 329.7833, 329.8633, 330.0033, 330.1433, 330.2833, 
    330.4333, 330.5833, 330.6733, 330.6933, 330.6833, 330.6833, 330.7333, 
    330.8633, 331.0633, 331.2633, 331.4633, 331.6633, 331.7833, 331.7433, 
    331.6633, 331.6133, 331.6333, 331.7233, 331.8433, 331.8833, 331.9233, 
    332.0733, 332.2633, 332.4133, 332.5092, 332.5692, 332.6292, 332.7092, 
    332.7792, 332.8892, 333.0292, 333.1592, 333.2592, 333.4192, 333.6192, 
    333.7892, 333.9075, 333.9875, 334.0375, 334.0875, 334.1275, 334.1475, 
    334.1675, 334.2575, 334.4275, 334.6375, 334.8575, 335.0775, 335.25, 
    335.35, 335.41, 335.46, 335.47, 335.49, 335.55, 335.64, 335.76, 335.93, 
    336.15, 336.34, 336.47, 336.53, 336.57, 336.58, 336.56, 336.58, 336.62,
    336.66, 336.73, 336.88, 337.09, 337.31 ;

 year = 1750.083, 1750.167, 1750.25, 1750.333, 1750.417, 1750.5, 1750.583, 
    1750.667, 1750.75, 1750.833, 1750.917, 1751, 1751.083, 1751.167, 1751.25, 
    1751.333, 1751.417, 1751.5, 1751.583, 1751.667, 1751.75, 1751.833, 
    1751.917, 1752, 1752.083, 1752.167, 1752.25, 1752.333, 1752.417, 1752.5, 
    1752.583, 1752.667, 1752.75, 1752.833, 1752.917, 1753, 1753.083, 
    1753.167, 1753.25, 1753.333, 1753.417, 1753.5, 1753.583, 1753.667, 
    1753.75, 1753.833, 1753.917, 1754, 1754.083, 1754.167, 1754.25, 1754.333, 
    1754.417, 1754.5, 1754.583, 1754.667, 1754.75, 1754.833, 1754.917, 1755, 
    1755.083, 1755.167, 1755.25, 1755.333, 1755.417, 1755.5, 1755.583, 
    1755.667, 1755.75, 1755.833, 1755.917, 1756, 1756.083, 1756.167, 1756.25, 
    1756.333, 1756.417, 1756.5, 1756.583, 1756.667, 1756.75, 1756.833, 
    1756.917, 1757, 1757.083, 1757.167, 1757.25, 1757.333, 1757.417, 1757.5, 
    1757.583, 1757.667, 1757.75, 1757.833, 1757.917, 1758, 1758.083, 
    1758.167, 1758.25, 1758.333, 1758.417, 1758.5, 1758.583, 1758.667, 
    1758.75, 1758.833, 1758.917, 1759, 1759.083, 1759.167, 1759.25, 1759.333, 
    1759.417, 1759.5, 1759.583, 1759.667, 1759.75, 1759.833, 1759.917, 1760, 
    1760.083, 1760.167, 1760.25, 1760.333, 1760.417, 1760.5, 1760.583, 
    1760.667, 1760.75, 1760.833, 1760.917, 1761, 1761.083, 1761.167, 1761.25, 
    1761.333, 1761.417, 1761.5, 1761.583, 1761.667, 1761.75, 1761.833, 
    1761.917, 1762, 1762.083, 1762.167, 1762.25, 1762.333, 1762.417, 1762.5, 
    1762.583, 1762.667, 1762.75, 1762.833, 1762.917, 1763, 1763.083, 
    1763.167, 1763.25, 1763.333, 1763.417, 1763.5, 1763.583, 1763.667, 
    1763.75, 1763.833, 1763.917, 1764, 1764.083, 1764.167, 1764.25, 1764.333, 
    1764.417, 1764.5, 1764.583, 1764.667, 1764.75, 1764.833, 1764.917, 1765, 
    1765.083, 1765.167, 1765.25, 1765.333, 1765.417, 1765.5, 1765.583, 
    1765.667, 1765.75, 1765.833, 1765.917, 1766, 1766.083, 1766.167, 1766.25, 
    1766.333, 1766.417, 1766.5, 1766.583, 1766.667, 1766.75, 1766.833, 
    1766.917, 1767, 1767.083, 1767.167, 1767.25, 1767.333, 1767.417, 1767.5, 
    1767.583, 1767.667, 1767.75, 1767.833, 1767.917, 1768, 1768.083, 
    1768.167, 1768.25, 1768.333, 1768.417, 1768.5, 1768.583, 1768.667, 
    1768.75, 1768.833, 1768.917, 1769, 1769.083, 1769.167, 1769.25, 1769.333, 
    1769.417, 1769.5, 1769.583, 1769.667, 1769.75, 1769.833, 1769.917, 1770, 
    1770.083, 1770.167, 1770.25, 1770.333, 1770.417, 1770.5, 1770.583, 
    1770.667, 1770.75, 1770.833, 1770.917, 1771, 1771.083, 1771.167, 1771.25, 
    1771.333, 1771.417, 1771.5, 1771.583, 1771.667, 1771.75, 1771.833, 
    1771.917, 1772, 1772.083, 1772.167, 1772.25, 1772.333, 1772.417, 1772.5, 
    1772.583, 1772.667, 1772.75, 1772.833, 1772.917, 1773, 1773.083, 
    1773.167, 1773.25, 1773.333, 1773.417, 1773.5, 1773.583, 1773.667, 
    1773.75, 1773.833, 1773.917, 1774, 1774.083, 1774.167, 1774.25, 1774.333, 
    1774.417, 1774.5, 1774.583, 1774.667, 1774.75, 1774.833, 1774.917, 1775, 
    1775.083, 1775.167, 1775.25, 1775.333, 1775.417, 1775.5, 1775.583, 
    1775.667, 1775.75, 1775.833, 1775.917, 1776, 1776.083, 1776.167, 1776.25, 
    1776.333, 1776.417, 1776.5, 1776.583, 1776.667, 1776.75, 1776.833, 
    1776.917, 1777, 1777.083, 1777.167, 1777.25, 1777.333, 1777.417, 1777.5, 
    1777.583, 1777.667, 1777.75, 1777.833, 1777.917, 1778, 1778.083, 
    1778.167, 1778.25, 1778.333, 1778.417, 1778.5, 1778.583, 1778.667, 
    1778.75, 1778.833, 1778.917, 1779, 1779.083, 1779.167, 1779.25, 1779.333, 
    1779.417, 1779.5, 1779.583, 1779.667, 1779.75, 1779.833, 1779.917, 1780, 
    1780.083, 1780.167, 1780.25, 1780.333, 1780.417, 1780.5, 1780.583, 
    1780.667, 1780.75, 1780.833, 1780.917, 1781, 1781.083, 1781.167, 1781.25, 
    1781.333, 1781.417, 1781.5, 1781.583, 1781.667, 1781.75, 1781.833, 
    1781.917, 1782, 1782.083, 1782.167, 1782.25, 1782.333, 1782.417, 1782.5, 
    1782.583, 1782.667, 1782.75, 1782.833, 1782.917, 1783, 1783.083, 
    1783.167, 1783.25, 1783.333, 1783.417, 1783.5, 1783.583, 1783.667, 
    1783.75, 1783.833, 1783.917, 1784, 1784.083, 1784.167, 1784.25, 1784.333, 
    1784.417, 1784.5, 1784.583, 1784.667, 1784.75, 1784.833, 1784.917, 1785, 
    1785.083, 1785.167, 1785.25, 1785.333, 1785.417, 1785.5, 1785.583, 
    1785.667, 1785.75, 1785.833, 1785.917, 1786, 1786.083, 1786.167, 1786.25, 
    1786.333, 1786.417, 1786.5, 1786.583, 1786.667, 1786.75, 1786.833, 
    1786.917, 1787, 1787.083, 1787.167, 1787.25, 1787.333, 1787.417, 1787.5, 
    1787.583, 1787.667, 1787.75, 1787.833, 1787.917, 1788, 1788.083, 
    1788.167, 1788.25, 1788.333, 1788.417, 1788.5, 1788.583, 1788.667, 
    1788.75, 1788.833, 1788.917, 1789, 1789.083, 1789.167, 1789.25, 1789.333, 
    1789.417, 1789.5, 1789.583, 1789.667, 1789.75, 1789.833, 1789.917, 1790, 
    1790.083, 1790.167, 1790.25, 1790.333, 1790.417, 1790.5, 1790.583, 
    1790.667, 1790.75, 1790.833, 1790.917, 1791, 1791.083, 1791.167, 1791.25, 
    1791.333, 1791.417, 1791.5, 1791.583, 1791.667, 1791.75, 1791.833, 
    1791.917, 1792, 1792.083, 1792.167, 1792.25, 1792.333, 1792.417, 1792.5, 
    1792.583, 1792.667, 1792.75, 1792.833, 1792.917, 1793, 1793.083, 
    1793.167, 1793.25, 1793.333, 1793.417, 1793.5, 1793.583, 1793.667, 
    1793.75, 1793.833, 1793.917, 1794, 1794.083, 1794.167, 1794.25, 1794.333, 
    1794.417, 1794.5, 1794.583, 1794.667, 1794.75, 1794.833, 1794.917, 1795, 
    1795.083, 1795.167, 1795.25, 1795.333, 1795.417, 1795.5, 1795.583, 
    1795.667, 1795.75, 1795.833, 1795.917, 1796, 1796.083, 1796.167, 1796.25, 
    1796.333, 1796.417, 1796.5, 1796.583, 1796.667, 1796.75, 1796.833, 
    1796.917, 1797, 1797.083, 1797.167, 1797.25, 1797.333, 1797.417, 1797.5, 
    1797.583, 1797.667, 1797.75, 1797.833, 1797.917, 1798, 1798.083, 
    1798.167, 1798.25, 1798.333, 1798.417, 1798.5, 1798.583, 1798.667, 
    1798.75, 1798.833, 1798.917, 1799, 1799.083, 1799.167, 1799.25, 1799.333, 
    1799.417, 1799.5, 1799.583, 1799.667, 1799.75, 1799.833, 1799.917, 1800, 
    1800.083, 1800.167, 1800.25, 1800.333, 1800.417, 1800.5, 1800.583, 
    1800.667, 1800.75, 1800.833, 1800.917, 1801, 1801.083, 1801.167, 1801.25, 
    1801.333, 1801.417, 1801.5, 1801.583, 1801.667, 1801.75, 1801.833, 
    1801.917, 1802, 1802.083, 1802.167, 1802.25, 1802.333, 1802.417, 1802.5, 
    1802.583, 1802.667, 1802.75, 1802.833, 1802.917, 1803, 1803.083, 
    1803.167, 1803.25, 1803.333, 1803.417, 1803.5, 1803.583, 1803.667, 
    1803.75, 1803.833, 1803.917, 1804, 1804.083, 1804.167, 1804.25, 1804.333, 
    1804.417, 1804.5, 1804.583, 1804.667, 1804.75, 1804.833, 1804.917, 1805, 
    1805.083, 1805.167, 1805.25, 1805.333, 1805.417, 1805.5, 1805.583, 
    1805.667, 1805.75, 1805.833, 1805.917, 1806, 1806.083, 1806.167, 1806.25, 
    1806.333, 1806.417, 1806.5, 1806.583, 1806.667, 1806.75, 1806.833, 
    1806.917, 1807, 1807.083, 1807.167, 1807.25, 1807.333, 1807.417, 1807.5, 
    1807.583, 1807.667, 1807.75, 1807.833, 1807.917, 1808, 1808.083, 
    1808.167, 1808.25, 1808.333, 1808.417, 1808.5, 1808.583, 1808.667, 
    1808.75, 1808.833, 1808.917, 1809, 1809.083, 1809.167, 1809.25, 1809.333, 
    1809.417, 1809.5, 1809.583, 1809.667, 1809.75, 1809.833, 1809.917, 1810, 
    1810.083, 1810.167, 1810.25, 1810.333, 1810.417, 1810.5, 1810.583, 
    1810.667, 1810.75, 1810.833, 1810.917, 1811, 1811.083, 1811.167, 1811.25, 
    1811.333, 1811.417, 1811.5, 1811.583, 1811.667, 1811.75, 1811.833, 
    1811.917, 1812, 1812.083, 1812.167, 1812.25, 1812.333, 1812.417, 1812.5, 
    1812.583, 1812.667, 1812.75, 1812.833, 1812.917, 1813, 1813.083, 
    1813.167, 1813.25, 1813.333, 1813.417, 1813.5, 1813.583, 1813.667, 
    1813.75, 1813.833, 1813.917, 1814, 1814.083, 1814.167, 1814.25, 1814.333, 
    1814.417, 1814.5, 1814.583, 1814.667, 1814.75, 1814.833, 1814.917, 1815, 
    1815.083, 1815.167, 1815.25, 1815.333, 1815.417, 1815.5, 1815.583, 
    1815.667, 1815.75, 1815.833, 1815.917, 1816, 1816.083, 1816.167, 1816.25, 
    1816.333, 1816.417, 1816.5, 1816.583, 1816.667, 1816.75, 1816.833, 
    1816.917, 1817, 1817.083, 1817.167, 1817.25, 1817.333, 1817.417, 1817.5, 
    1817.583, 1817.667, 1817.75, 1817.833, 1817.917, 1818, 1818.083, 
    1818.167, 1818.25, 1818.333, 1818.417, 1818.5, 1818.583, 1818.667, 
    1818.75, 1818.833, 1818.917, 1819, 1819.083, 1819.167, 1819.25, 1819.333, 
    1819.417, 1819.5, 1819.583, 1819.667, 1819.75, 1819.833, 1819.917, 1820, 
    1820.083, 1820.167, 1820.25, 1820.333, 1820.417, 1820.5, 1820.583, 
    1820.667, 1820.75, 1820.833, 1820.917, 1821, 1821.083, 1821.167, 1821.25, 
    1821.333, 1821.417, 1821.5, 1821.583, 1821.667, 1821.75, 1821.833, 
    1821.917, 1822, 1822.083, 1822.167, 1822.25, 1822.333, 1822.417, 1822.5, 
    1822.583, 1822.667, 1822.75, 1822.833, 1822.917, 1823, 1823.083, 
    1823.167, 1823.25, 1823.333, 1823.417, 1823.5, 1823.583, 1823.667, 
    1823.75, 1823.833, 1823.917, 1824, 1824.083, 1824.167, 1824.25, 1824.333, 
    1824.417, 1824.5, 1824.583, 1824.667, 1824.75, 1824.833, 1824.917, 1825, 
    1825.083, 1825.167, 1825.25, 1825.333, 1825.417, 1825.5, 1825.583, 
    1825.667, 1825.75, 1825.833, 1825.917, 1826, 1826.083, 1826.167, 1826.25, 
    1826.333, 1826.417, 1826.5, 1826.583, 1826.667, 1826.75, 1826.833, 
    1826.917, 1827, 1827.083, 1827.167, 1827.25, 1827.333, 1827.417, 1827.5, 
    1827.583, 1827.667, 1827.75, 1827.833, 1827.917, 1828, 1828.083, 
    1828.167, 1828.25, 1828.333, 1828.417, 1828.5, 1828.583, 1828.667, 
    1828.75, 1828.833, 1828.917, 1829, 1829.083, 1829.167, 1829.25, 1829.333, 
    1829.417, 1829.5, 1829.583, 1829.667, 1829.75, 1829.833, 1829.917, 1830, 
    1830.083, 1830.167, 1830.25, 1830.333, 1830.417, 1830.5, 1830.583, 
    1830.667, 1830.75, 1830.833, 1830.917, 1831, 1831.083, 1831.167, 1831.25, 
    1831.333, 1831.417, 1831.5, 1831.583, 1831.667, 1831.75, 1831.833, 
    1831.917, 1832, 1832.083, 1832.167, 1832.25, 1832.333, 1832.417, 1832.5, 
    1832.583, 1832.667, 1832.75, 1832.833, 1832.917, 1833, 1833.083, 
    1833.167, 1833.25, 1833.333, 1833.417, 1833.5, 1833.583, 1833.667, 
    1833.75, 1833.833, 1833.917, 1834, 1834.083, 1834.167, 1834.25, 1834.333, 
    1834.417, 1834.5, 1834.583, 1834.667, 1834.75, 1834.833, 1834.917, 1835, 
    1835.083, 1835.167, 1835.25, 1835.333, 1835.417, 1835.5, 1835.583, 
    1835.667, 1835.75, 1835.833, 1835.917, 1836, 1836.083, 1836.167, 1836.25, 
    1836.333, 1836.417, 1836.5, 1836.583, 1836.667, 1836.75, 1836.833, 
    1836.917, 1837, 1837.083, 1837.167, 1837.25, 1837.333, 1837.417, 1837.5, 
    1837.583, 1837.667, 1837.75, 1837.833, 1837.917, 1838, 1838.083, 
    1838.167, 1838.25, 1838.333, 1838.417, 1838.5, 1838.583, 1838.667, 
    1838.75, 1838.833, 1838.917, 1839, 1839.083, 1839.167, 1839.25, 1839.333, 
    1839.417, 1839.5, 1839.583, 1839.667, 1839.75, 1839.833, 1839.917, 1840, 
    1840.083, 1840.167, 1840.25, 1840.333, 1840.417, 1840.5, 1840.583, 
    1840.667, 1840.75, 1840.833, 1840.917, 1841, 1841.083, 1841.167, 1841.25, 
    1841.333, 1841.417, 1841.5, 1841.583, 1841.667, 1841.75, 1841.833, 
    1841.917, 1842, 1842.083, 1842.167, 1842.25, 1842.333, 1842.417, 1842.5, 
    1842.583, 1842.667, 1842.75, 1842.833, 1842.917, 1843, 1843.083, 
    1843.167, 1843.25, 1843.333, 1843.417, 1843.5, 1843.583, 1843.667, 
    1843.75, 1843.833, 1843.917, 1844, 1844.083, 1844.167, 1844.25, 1844.333, 
    1844.417, 1844.5, 1844.583, 1844.667, 1844.75, 1844.833, 1844.917, 1845, 
    1845.083, 1845.167, 1845.25, 1845.333, 1845.417, 1845.5, 1845.583, 
    1845.667, 1845.75, 1845.833, 1845.917, 1846, 1846.083, 1846.167, 1846.25, 
    1846.333, 1846.417, 1846.5, 1846.583, 1846.667, 1846.75, 1846.833, 
    1846.917, 1847, 1847.083, 1847.167, 1847.25, 1847.333, 1847.417, 1847.5, 
    1847.583, 1847.667, 1847.75, 1847.833, 1847.917, 1848, 1848.083, 
    1848.167, 1848.25, 1848.333, 1848.417, 1848.5, 1848.583, 1848.667, 
    1848.75, 1848.833, 1848.917, 1849, 1849.083, 1849.167, 1849.25, 1849.333, 
    1849.417, 1849.5, 1849.583, 1849.667, 1849.75, 1849.833, 1849.917, 1850, 
    1850.083, 1850.167, 1850.25, 1850.333, 1850.417, 1850.5, 1850.583, 
    1850.667, 1850.75, 1850.833, 1850.917, 1851, 1851.083, 1851.167, 1851.25, 
    1851.333, 1851.417, 1851.5, 1851.583, 1851.667, 1851.75, 1851.833, 
    1851.917, 1852, 1852.083, 1852.167, 1852.25, 1852.333, 1852.417, 1852.5, 
    1852.583, 1852.667, 1852.75, 1852.833, 1852.917, 1853, 1853.083, 
    1853.167, 1853.25, 1853.333, 1853.417, 1853.5, 1853.583, 1853.667, 
    1853.75, 1853.833, 1853.917, 1854, 1854.083, 1854.167, 1854.25, 1854.333, 
    1854.417, 1854.5, 1854.583, 1854.667, 1854.75, 1854.833, 1854.917, 1855, 
    1855.083, 1855.167, 1855.25, 1855.333, 1855.417, 1855.5, 1855.583, 
    1855.667, 1855.75, 1855.833, 1855.917, 1856, 1856.083, 1856.167, 1856.25, 
    1856.333, 1856.417, 1856.5, 1856.583, 1856.667, 1856.75, 1856.833, 
    1856.917, 1857, 1857.083, 1857.167, 1857.25, 1857.333, 1857.417, 1857.5, 
    1857.583, 1857.667, 1857.75, 1857.833, 1857.917, 1858, 1858.083, 
    1858.167, 1858.25, 1858.333, 1858.417, 1858.5, 1858.583, 1858.667, 
    1858.75, 1858.833, 1858.917, 1859, 1859.083, 1859.167, 1859.25, 1859.333, 
    1859.417, 1859.5, 1859.583, 1859.667, 1859.75, 1859.833, 1859.917, 1860, 
    1860.083, 1860.167, 1860.25, 1860.333, 1860.417, 1860.5, 1860.583, 
    1860.667, 1860.75, 1860.833, 1860.917, 1861, 1861.083, 1861.167, 1861.25, 
    1861.333, 1861.417, 1861.5, 1861.583, 1861.667, 1861.75, 1861.833, 
    1861.917, 1862, 1862.083, 1862.167, 1862.25, 1862.333, 1862.417, 1862.5, 
    1862.583, 1862.667, 1862.75, 1862.833, 1862.917, 1863, 1863.083, 
    1863.167, 1863.25, 1863.333, 1863.417, 1863.5, 1863.583, 1863.667, 
    1863.75, 1863.833, 1863.917, 1864, 1864.083, 1864.167, 1864.25, 1864.333, 
    1864.417, 1864.5, 1864.583, 1864.667, 1864.75, 1864.833, 1864.917, 1865, 
    1865.083, 1865.167, 1865.25, 1865.333, 1865.417, 1865.5, 1865.583, 
    1865.667, 1865.75, 1865.833, 1865.917, 1866, 1866.083, 1866.167, 1866.25, 
    1866.333, 1866.417, 1866.5, 1866.583, 1866.667, 1866.75, 1866.833, 
    1866.917, 1867, 1867.083, 1867.167, 1867.25, 1867.333, 1867.417, 1867.5, 
    1867.583, 1867.667, 1867.75, 1867.833, 1867.917, 1868, 1868.083, 
    1868.167, 1868.25, 1868.333, 1868.417, 1868.5, 1868.583, 1868.667, 
    1868.75, 1868.833, 1868.917, 1869, 1869.083, 1869.167, 1869.25, 1869.333, 
    1869.417, 1869.5, 1869.583, 1869.667, 1869.75, 1869.833, 1869.917, 1870, 
    1870.083, 1870.167, 1870.25, 1870.333, 1870.417, 1870.5, 1870.583, 
    1870.667, 1870.75, 1870.833, 1870.917, 1871, 1871.083, 1871.167, 1871.25, 
    1871.333, 1871.417, 1871.5, 1871.583, 1871.667, 1871.75, 1871.833, 
    1871.917, 1872, 1872.083, 1872.167, 1872.25, 1872.333, 1872.417, 1872.5, 
    1872.583, 1872.667, 1872.75, 1872.833, 1872.917, 1873, 1873.083, 
    1873.167, 1873.25, 1873.333, 1873.417, 1873.5, 1873.583, 1873.667, 
    1873.75, 1873.833, 1873.917, 1874, 1874.083, 1874.167, 1874.25, 1874.333, 
    1874.417, 1874.5, 1874.583, 1874.667, 1874.75, 1874.833, 1874.917, 1875, 
    1875.083, 1875.167, 1875.25, 1875.333, 1875.417, 1875.5, 1875.583, 
    1875.667, 1875.75, 1875.833, 1875.917, 1876, 1876.083, 1876.167, 1876.25, 
    1876.333, 1876.417, 1876.5, 1876.583, 1876.667, 1876.75, 1876.833, 
    1876.917, 1877, 1877.083, 1877.167, 1877.25, 1877.333, 1877.417, 1877.5, 
    1877.583, 1877.667, 1877.75, 1877.833, 1877.917, 1878, 1878.083, 
    1878.167, 1878.25, 1878.333, 1878.417, 1878.5, 1878.583, 1878.667, 
    1878.75, 1878.833, 1878.917, 1879, 1879.083, 1879.167, 1879.25, 1879.333, 
    1879.417, 1879.5, 1879.583, 1879.667, 1879.75, 1879.833, 1879.917, 1880, 
    1880.083, 1880.167, 1880.25, 1880.333, 1880.417, 1880.5, 1880.583, 
    1880.667, 1880.75, 1880.833, 1880.917, 1881, 1881.083, 1881.167, 1881.25, 
    1881.333, 1881.417, 1881.5, 1881.583, 1881.667, 1881.75, 1881.833, 
    1881.917, 1882, 1882.083, 1882.167, 1882.25, 1882.333, 1882.417, 1882.5, 
    1882.583, 1882.667, 1882.75, 1882.833, 1882.917, 1883, 1883.083, 
    1883.167, 1883.25, 1883.333, 1883.417, 1883.5, 1883.583, 1883.667, 
    1883.75, 1883.833, 1883.917, 1884, 1884.083, 1884.167, 1884.25, 1884.333, 
    1884.417, 1884.5, 1884.583, 1884.667, 1884.75, 1884.833, 1884.917, 1885, 
    1885.083, 1885.167, 1885.25, 1885.333, 1885.417, 1885.5, 1885.583, 
    1885.667, 1885.75, 1885.833, 1885.917, 1886, 1886.083, 1886.167, 1886.25, 
    1886.333, 1886.417, 1886.5, 1886.583, 1886.667, 1886.75, 1886.833, 
    1886.917, 1887, 1887.083, 1887.167, 1887.25, 1887.333, 1887.417, 1887.5, 
    1887.583, 1887.667, 1887.75, 1887.833, 1887.917, 1888, 1888.083, 
    1888.167, 1888.25, 1888.333, 1888.417, 1888.5, 1888.583, 1888.667, 
    1888.75, 1888.833, 1888.917, 1889, 1889.083, 1889.167, 1889.25, 1889.333, 
    1889.417, 1889.5, 1889.583, 1889.667, 1889.75, 1889.833, 1889.917, 1890, 
    1890.083, 1890.167, 1890.25, 1890.333, 1890.417, 1890.5, 1890.583, 
    1890.667, 1890.75, 1890.833, 1890.917, 1891, 1891.083, 1891.167, 1891.25, 
    1891.333, 1891.417, 1891.5, 1891.583, 1891.667, 1891.75, 1891.833, 
    1891.917, 1892, 1892.083, 1892.167, 1892.25, 1892.333, 1892.417, 1892.5, 
    1892.583, 1892.667, 1892.75, 1892.833, 1892.917, 1893, 1893.083, 
    1893.167, 1893.25, 1893.333, 1893.417, 1893.5, 1893.583, 1893.667, 
    1893.75, 1893.833, 1893.917, 1894, 1894.083, 1894.167, 1894.25, 1894.333, 
    1894.417, 1894.5, 1894.583, 1894.667, 1894.75, 1894.833, 1894.917, 1895, 
    1895.083, 1895.167, 1895.25, 1895.333, 1895.417, 1895.5, 1895.583, 
    1895.667, 1895.75, 1895.833, 1895.917, 1896, 1896.083, 1896.167, 1896.25, 
    1896.333, 1896.417, 1896.5, 1896.583, 1896.667, 1896.75, 1896.833, 
    1896.917, 1897, 1897.083, 1897.167, 1897.25, 1897.333, 1897.417, 1897.5, 
    1897.583, 1897.667, 1897.75, 1897.833, 1897.917, 1898, 1898.083, 
    1898.167, 1898.25, 1898.333, 1898.417, 1898.5, 1898.583, 1898.667, 
    1898.75, 1898.833, 1898.917, 1899, 1899.083, 1899.167, 1899.25, 1899.333, 
    1899.417, 1899.5, 1899.583, 1899.667, 1899.75, 1899.833, 1899.917, 1900, 
    1900.083, 1900.167, 1900.25, 1900.333, 1900.417, 1900.5, 1900.583, 
    1900.667, 1900.75, 1900.833, 1900.917, 1901, 1901.083, 1901.167, 1901.25, 
    1901.333, 1901.417, 1901.5, 1901.583, 1901.667, 1901.75, 1901.833, 
    1901.917, 1902, 1902.083, 1902.167, 1902.25, 1902.333, 1902.417, 1902.5, 
    1902.583, 1902.667, 1902.75, 1902.833, 1902.917, 1903, 1903.083, 
    1903.167, 1903.25, 1903.333, 1903.417, 1903.5, 1903.583, 1903.667, 
    1903.75, 1903.833, 1903.917, 1904, 1904.083, 1904.167, 1904.25, 1904.333, 
    1904.417, 1904.5, 1904.583, 1904.667, 1904.75, 1904.833, 1904.917, 1905, 
    1905.083, 1905.167, 1905.25, 1905.333, 1905.417, 1905.5, 1905.583, 
    1905.667, 1905.75, 1905.833, 1905.917, 1906, 1906.083, 1906.167, 1906.25, 
    1906.333, 1906.417, 1906.5, 1906.583, 1906.667, 1906.75, 1906.833, 
    1906.917, 1907, 1907.083, 1907.167, 1907.25, 1907.333, 1907.417, 1907.5, 
    1907.583, 1907.667, 1907.75, 1907.833, 1907.917, 1908, 1908.083, 
    1908.167, 1908.25, 1908.333, 1908.417, 1908.5, 1908.583, 1908.667, 
    1908.75, 1908.833, 1908.917, 1909, 1909.083, 1909.167, 1909.25, 1909.333, 
    1909.417, 1909.5, 1909.583, 1909.667, 1909.75, 1909.833, 1909.917, 1910, 
    1910.083, 1910.167, 1910.25, 1910.333, 1910.417, 1910.5, 1910.583, 
    1910.667, 1910.75, 1910.833, 1910.917, 1911, 1911.083, 1911.167, 1911.25, 
    1911.333, 1911.417, 1911.5, 1911.583, 1911.667, 1911.75, 1911.833, 
    1911.917, 1912, 1912.083, 1912.167, 1912.25, 1912.333, 1912.417, 1912.5, 
    1912.583, 1912.667, 1912.75, 1912.833, 1912.917, 1913, 1913.083, 
    1913.167, 1913.25, 1913.333, 1913.417, 1913.5, 1913.583, 1913.667, 
    1913.75, 1913.833, 1913.917, 1914, 1914.083, 1914.167, 1914.25, 1914.333, 
    1914.417, 1914.5, 1914.583, 1914.667, 1914.75, 1914.833, 1914.917, 1915, 
    1915.083, 1915.167, 1915.25, 1915.333, 1915.417, 1915.5, 1915.583, 
    1915.667, 1915.75, 1915.833, 1915.917, 1916, 1916.083, 1916.167, 1916.25, 
    1916.333, 1916.417, 1916.5, 1916.583, 1916.667, 1916.75, 1916.833, 
    1916.917, 1917, 1917.083, 1917.167, 1917.25, 1917.333, 1917.417, 1917.5, 
    1917.583, 1917.667, 1917.75, 1917.833, 1917.917, 1918, 1918.083, 
    1918.167, 1918.25, 1918.333, 1918.417, 1918.5, 1918.583, 1918.667, 
    1918.75, 1918.833, 1918.917, 1919, 1919.083, 1919.167, 1919.25, 1919.333, 
    1919.417, 1919.5, 1919.583, 1919.667, 1919.75, 1919.833, 1919.917, 1920, 
    1920.083, 1920.167, 1920.25, 1920.333, 1920.417, 1920.5, 1920.583, 
    1920.667, 1920.75, 1920.833, 1920.917, 1921, 1921.083, 1921.167, 1921.25, 
    1921.333, 1921.417, 1921.5, 1921.583, 1921.667, 1921.75, 1921.833, 
    1921.917, 1922, 1922.083, 1922.167, 1922.25, 1922.333, 1922.417, 1922.5, 
    1922.583, 1922.667, 1922.75, 1922.833, 1922.917, 1923, 1923.083, 
    1923.167, 1923.25, 1923.333, 1923.417, 1923.5, 1923.583, 1923.667, 
    1923.75, 1923.833, 1923.917, 1924, 1924.083, 1924.167, 1924.25, 1924.333, 
    1924.417, 1924.5, 1924.583, 1924.667, 1924.75, 1924.833, 1924.917, 1925, 
    1925.083, 1925.167, 1925.25, 1925.333, 1925.417, 1925.5, 1925.583, 
    1925.667, 1925.75, 1925.833, 1925.917, 1926, 1926.083, 1926.167, 1926.25, 
    1926.333, 1926.417, 1926.5, 1926.583, 1926.667, 1926.75, 1926.833, 
    1926.917, 1927, 1927.083, 1927.167, 1927.25, 1927.333, 1927.417, 1927.5, 
    1927.583, 1927.667, 1927.75, 1927.833, 1927.917, 1928, 1928.083, 
    1928.167, 1928.25, 1928.333, 1928.417, 1928.5, 1928.583, 1928.667, 
    1928.75, 1928.833, 1928.917, 1929, 1929.083, 1929.167, 1929.25, 1929.333, 
    1929.417, 1929.5, 1929.583, 1929.667, 1929.75, 1929.833, 1929.917, 1930, 
    1930.083, 1930.167, 1930.25, 1930.333, 1930.417, 1930.5, 1930.583, 
    1930.667, 1930.75, 1930.833, 1930.917, 1931, 1931.083, 1931.167, 1931.25, 
    1931.333, 1931.417, 1931.5, 1931.583, 1931.667, 1931.75, 1931.833, 
    1931.917, 1932, 1932.083, 1932.167, 1932.25, 1932.333, 1932.417, 1932.5, 
    1932.583, 1932.667, 1932.75, 1932.833, 1932.917, 1933, 1933.083, 
    1933.167, 1933.25, 1933.333, 1933.417, 1933.5, 1933.583, 1933.667, 
    1933.75, 1933.833, 1933.917, 1934, 1934.083, 1934.167, 1934.25, 1934.333, 
    1934.417, 1934.5, 1934.583, 1934.667, 1934.75, 1934.833, 1934.917, 1935, 
    1935.083, 1935.167, 1935.25, 1935.333, 1935.417, 1935.5, 1935.583, 
    1935.667, 1935.75, 1935.833, 1935.917, 1936, 1936.083, 1936.167, 1936.25, 
    1936.333, 1936.417, 1936.5, 1936.583, 1936.667, 1936.75, 1936.833, 
    1936.917, 1937, 1937.083, 1937.167, 1937.25, 1937.333, 1937.417, 1937.5, 
    1937.583, 1937.667, 1937.75, 1937.833, 1937.917, 1938, 1938.083, 
    1938.167, 1938.25, 1938.333, 1938.417, 1938.5, 1938.583, 1938.667, 
    1938.75, 1938.833, 1938.917, 1939, 1939.083, 1939.167, 1939.25, 1939.333, 
    1939.417, 1939.5, 1939.583, 1939.667, 1939.75, 1939.833, 1939.917, 1940, 
    1940.083, 1940.167, 1940.25, 1940.333, 1940.417, 1940.5, 1940.583, 
    1940.667, 1940.75, 1940.833, 1940.917, 1941, 1941.083, 1941.167, 1941.25, 
    1941.333, 1941.417, 1941.5, 1941.583, 1941.667, 1941.75, 1941.833, 
    1941.917, 1942, 1942.083, 1942.167, 1942.25, 1942.333, 1942.417, 1942.5, 
    1942.583, 1942.667, 1942.75, 1942.833, 1942.917, 1943, 1943.083, 
    1943.167, 1943.25, 1943.333, 1943.417, 1943.5, 1943.583, 1943.667, 
    1943.75, 1943.833, 1943.917, 1944, 1944.083, 1944.167, 1944.25, 1944.333, 
    1944.417, 1944.5, 1944.583, 1944.667, 1944.75, 1944.833, 1944.917, 1945, 
    1945.083, 1945.167, 1945.25, 1945.333, 1945.417, 1945.5, 1945.583, 
    1945.667, 1945.75, 1945.833, 1945.917, 1946, 1946.083, 1946.167, 1946.25, 
    1946.333, 1946.417, 1946.5, 1946.583, 1946.667, 1946.75, 1946.833, 
    1946.917, 1947, 1947.083, 1947.167, 1947.25, 1947.333, 1947.417, 1947.5, 
    1947.583, 1947.667, 1947.75, 1947.833, 1947.917, 1948, 1948.083, 
    1948.167, 1948.25, 1948.333, 1948.417, 1948.5, 1948.583, 1948.667, 
    1948.75, 1948.833, 1948.917, 1949, 1949.083, 1949.167, 1949.25, 1949.333, 
    1949.417, 1949.5, 1949.583, 1949.667, 1949.75, 1949.833, 1949.917, 1950, 
    1950.083, 1950.167, 1950.25, 1950.333, 1950.417, 1950.5, 1950.583, 
    1950.667, 1950.75, 1950.833, 1950.917, 1951, 1951.083, 1951.167, 1951.25, 
    1951.333, 1951.417, 1951.5, 1951.583, 1951.667, 1951.75, 1951.833, 
    1951.917, 1952, 1952.083, 1952.167, 1952.25, 1952.333, 1952.417, 1952.5, 
    1952.583, 1952.667, 1952.75, 1952.833, 1952.917, 1953, 1953.083, 
    1953.167, 1953.25, 1953.333, 1953.417, 1953.5, 1953.583, 1953.667, 
    1953.75, 1953.833, 1953.917, 1954, 1954.083, 1954.167, 1954.25, 1954.333, 
    1954.417, 1954.5, 1954.583, 1954.667, 1954.75, 1954.833, 1954.917, 1955, 
    1955.083, 1955.167, 1955.25, 1955.333, 1955.417, 1955.5, 1955.583, 
    1955.667, 1955.75, 1955.833, 1955.917, 1956, 1956.083, 1956.167, 1956.25, 
    1956.333, 1956.417, 1956.5, 1956.583, 1956.667, 1956.75, 1956.833, 
    1956.917, 1957, 1957.083, 1957.167, 1957.25, 1957.333, 1957.417, 1957.5, 
    1957.583, 1957.667, 1957.75, 1957.833, 1957.917, 1958, 1958.083, 
    1958.167, 1958.25, 1958.333, 1958.417, 1958.5, 1958.583, 1958.667, 
    1958.75, 1958.833, 1958.917, 1959, 1959.083, 1959.167, 1959.25, 1959.333, 
    1959.417, 1959.5, 1959.583, 1959.667, 1959.75, 1959.833, 1959.917, 1960, 
    1960.083, 1960.167, 1960.25, 1960.333, 1960.417, 1960.5, 1960.583, 
    1960.667, 1960.75, 1960.833, 1960.917, 1961, 1961.083, 1961.167, 1961.25, 
    1961.333, 1961.417, 1961.5, 1961.583, 1961.667, 1961.75, 1961.833, 
    1961.917, 1962, 1962.083, 1962.167, 1962.25, 1962.333, 1962.417, 1962.5, 
    1962.583, 1962.667, 1962.75, 1962.833, 1962.917, 1963, 1963.083, 
    1963.167, 1963.25, 1963.333, 1963.417, 1963.5, 1963.583, 1963.667, 
    1963.75, 1963.833, 1963.917, 1964, 1964.083, 1964.167, 1964.25, 1964.333, 
    1964.417, 1964.5, 1964.583, 1964.667, 1964.75, 1964.833, 1964.917, 1965, 
    1965.083, 1965.167, 1965.25, 1965.333, 1965.417, 1965.5, 1965.583, 
    1965.667, 1965.75, 1965.833, 1965.917, 1966, 1966.083, 1966.167, 1966.25, 
    1966.333, 1966.417, 1966.5, 1966.583, 1966.667, 1966.75, 1966.833, 
    1966.917, 1967, 1967.083, 1967.167, 1967.25, 1967.333, 1967.417, 1967.5, 
    1967.583, 1967.667, 1967.75, 1967.833, 1967.917, 1968, 1968.083, 
    1968.167, 1968.25, 1968.333, 1968.417, 1968.5, 1968.583, 1968.667, 
    1968.75, 1968.833, 1968.917, 1969, 1969.083, 1969.167, 1969.25, 1969.333, 
    1969.417, 1969.5, 1969.583, 1969.667, 1969.75, 1969.833, 1969.917, 1970, 
    1970.083, 1970.167, 1970.25, 1970.333, 1970.417, 1970.5, 1970.583, 
    1970.667, 1970.75, 1970.833, 1970.917, 1971, 1971.083, 1971.167, 1971.25, 
    1971.333, 1971.417, 1971.5, 1971.583, 1971.667, 1971.75, 1971.833, 
    1971.917, 1972, 1972.083, 1972.167, 1972.25, 1972.333, 1972.417, 1972.5, 
    1972.583, 1972.667, 1972.75, 1972.833, 1972.917, 1973, 1973.083, 
    1973.167, 1973.25, 1973.333, 1973.417, 1973.5, 1973.583, 1973.667, 
    1973.75, 1973.833, 1973.917, 1974, 1974.083, 1974.167, 1974.25, 1974.333, 
    1974.417, 1974.5, 1974.583, 1974.667, 1974.75, 1974.833, 1974.917, 1975, 
    1975.083, 1975.167, 1975.25, 1975.333, 1975.417, 1975.5, 1975.583, 
    1975.667, 1975.75, 1975.833, 1975.917, 1976, 1976.083, 1976.167, 1976.25, 
    1976.333, 1976.417, 1976.5, 1976.583, 1976.667, 1976.75, 1976.833, 
    1976.917, 1977, 1977.083, 1977.167, 1977.25, 1977.333, 1977.417, 1977.5, 
    1977.583, 1977.667, 1977.75, 1977.833, 1977.917, 1978, 1978.083, 
    1978.167, 1978.25, 1978.333, 1978.417, 1978.5, 1978.583, 1978.667, 
    1978.75, 1978.833, 1978.917, 1979, 1979.083, 1979.167, 1979.25, 1979.333, 
    1979.417, 1979.5, 1979.583, 1979.667, 1979.75, 1979.833, 1979.917, 1980, 
    1980.083, 1980.167, 1980.25, 1980.333, 1980.417, 1980.5, 1980.583, 
    1980.667, 1980.75, 1980.833, 1980.917, 1981, 1981.083, 1981.167, 1981.25, 
    1981.333, 1981.417, 1981.5, 1981.583, 1981.667, 1981.75, 1981.833, 
    1981.917, 1982, 1982.083, 1982.167, 1982.25, 1982.333, 1982.417, 1982.5, 
    1982.583, 1982.667, 1982.75, 1982.833, 1982.917, 1983, 1983.083, 
    1983.167, 1983.25, 1983.333, 1983.417, 1983.5, 1983.583, 1983.667, 
    1983.75, 1983.833, 1983.917, 1984, 1984.083, 1984.167, 1984.25, 1984.333, 
    1984.417, 1984.5, 1984.583, 1984.667, 1984.75, 1984.833, 1984.917, 1985, 
    1985.083, 1985.167, 1985.25, 1985.333, 1985.417, 1985.5, 1985.583, 
    1985.667, 1985.75, 1985.833, 1985.917, 1986, 1986.083, 1986.167, 1986.25, 
    1986.333, 1986.417, 1986.5, 1986.583, 1986.667, 1986.75, 1986.833, 
    1986.917, 1987, 1987.083, 1987.167, 1987.25, 1987.333, 1987.417, 1987.5, 
    1987.583, 1987.667, 1987.75, 1987.833, 1987.917, 1988, 1988.083, 
    1988.167, 1988.25, 1988.333, 1988.417, 1988.5, 1988.583, 1988.667, 
    1988.75, 1988.833, 1988.917, 1989, 1989.083, 1989.167, 1989.25, 1989.333, 
    1989.417, 1989.5, 1989.583, 1989.667, 1989.75, 1989.833, 1989.917, 1990, 
    1990.083, 1990.167, 1990.25, 1990.333, 1990.417, 1990.5, 1990.583, 
    1990.667, 1990.75, 1990.833, 1990.917, 1991, 1991.083, 1991.167, 1991.25, 
    1991.333, 1991.417, 1991.5, 1991.583, 1991.667, 1991.75, 1991.833, 
    1991.917, 1992, 1992.083, 1992.167, 1992.25, 1992.333, 1992.417, 1992.5, 
    1992.583, 1992.667, 1992.75, 1992.833, 1992.917, 1993, 1993.083, 
    1993.167, 1993.25, 1993.333, 1993.417, 1993.5, 1993.583, 1993.667, 
    1993.75, 1993.833, 1993.917, 1994, 1994.083, 1994.167, 1994.25, 1994.333, 
    1994.417, 1994.5, 1994.583, 1994.667, 1994.75, 1994.833, 1994.917, 1995, 
    1995.083, 1995.167, 1995.25, 1995.333, 1995.417, 1995.5, 1995.583, 
    1995.667, 1995.75, 1995.833, 1995.917, 1996, 1996.083, 1996.167, 1996.25, 
    1996.333, 1996.417, 1996.5, 1996.583, 1996.667, 1996.75, 1996.833, 
    1996.917, 1997, 1997.083, 1997.167, 1997.25, 1997.333, 1997.417, 1997.5, 
    1997.583, 1997.667, 1997.75, 1997.833, 1997.917, 1998, 1998.083, 
    1998.167, 1998.25, 1998.333, 1998.417, 1998.5, 1998.583, 1998.667, 
    1998.75, 1998.833, 1998.917, 1999, 1999.083, 1999.167, 1999.25, 1999.333, 
    1999.417, 1999.5, 1999.583, 1999.667, 1999.75, 1999.833, 1999.917, 2000, 
    2000.083, 2000.167, 2000.25, 2000.333, 2000.417, 2000.5, 2000.583, 
    2000.667, 2000.75, 2000.833, 2000.917, 2001, 2001.083, 2001.167, 2001.25, 
    2001.333, 2001.417, 2001.5, 2001.583, 2001.667, 2001.75, 2001.833, 
    2001.917, 2002, 2002.083, 2002.167, 2002.25, 2002.333, 2002.417, 2002.5, 
    2002.583, 2002.667, 2002.75, 2002.833, 2002.917, 2003, 2003.083, 
    2003.167, 2003.25, 2003.333, 2003.417, 2003.5, 2003.583, 2003.667, 
    2003.75, 2003.833, 2003.917, 2004, 2004.083, 2004.167, 2004.25, 2004.333, 
    2004.417, 2004.5, 2004.583, 2004.667, 2004.75, 2004.833, 2004.917, 2005, 
    2005.083, 2005.167, 2005.25, 2005.333, 2005.417, 2005.5, 2005.583, 
    2005.667, 2005.75, 2005.833, 2005.917, 2006, 2006.083, 2006.167, 2006.25, 
    2006.333, 2006.417, 2006.5, 2006.583, 2006.667, 2006.75, 2006.833, 
    2006.917, 2007, 2007.083, 2007.167, 2007.25, 2007.333, 2007.417, 2007.5, 
    2007.583, 2007.667, 2007.75, 2007.833, 2007.917, 2008, 2008.083, 
    2008.167, 2008.25, 2008.333, 2008.417, 2008.5, 2008.583, 2008.667, 
    2008.75, 2008.833, 2008.917, 2009, 2009.083, 2009.167, 2009.25, 2009.333, 
    2009.417, 2009.5, 2009.583, 2009.667, 2009.75, 2009.833, 2009.917, 2010, 
    2010.083, 2010.167, 2010.25, 2010.333, 2010.417, 2010.5, 2010.583, 
    2010.667, 2010.75, 2010.833, 2010.917, 2011, 2011.083, 2011.167, 2011.25, 
    2011.333, 2011.417, 2011.5, 2011.583, 2011.667, 2011.75, 2011.833, 
    2011.917, 2012, 2012.083, 2012.167, 2012.25, 2012.333, 2012.417, 2012.5, 
    2012.583, 2012.667, 2012.75, 2012.833, 2012.917, 2013, 2013.083, 
    2013.167, 2013.25, 2013.333, 2013.417, 2013.5, 2013.583, 2013.667, 
    2013.75, 2013.833, 2013.917, 2014, 2014.083, 2014.167, 2014.25, 2014.333, 
    2014.417, 2014.5, 2014.583, 2014.667, 2014.75, 2014.833, 2014.917, 2015, 
    2015.083, 2015.167, 2015.25, 2015.333, 2015.417, 2015.5, 2015.583, 
    2015.667, 2015.75, 2015.833, 2015.917, 2016, 2016.083, 2016.167, 2016.25, 
    2016.333, 2016.417, 2016.5, 2016.583, 2016.667, 2016.75, 2016.833, 
    2016.917, 2017, 2017.083, 2017.167, 2017.25, 2017.333, 2017.417, 2017.5, 
    2017.583, 2017.667, 2017.75, 2017.833, 2017.917, 2018, 2018.083, 
    2018.167, 2018.25, 2018.333, 2018.417, 2018.5, 2018.583, 2018.667, 
    2018.75, 2018.833, 2018.917, 2019, 2019.083, 2019.167, 2019.25, 2019.333, 
    2019.417, 2019.5, 2019.583, 2019.667, 2019.75, 2019.833, 2019.917, 2020, 
    2020.083, 2020.167, 2020.25, 2020.333, 2020.417, 2020.5, 2020.583, 
    2020.667, 2020.75, 2020.833, 2020.917, 2021, 2021.083, 2021.167, 2021.25, 
    2021.333, 2021.417, 2021.5, 2021.583, 2021.667, 2021.75, 2021.833, 
    2021.917, 2022, 2022.083, 2022.167, 2022.25, 2022.333, 2022.417, 2022.5, 
    2022.583, 2022.667, 2022.75, 2022.833, 2022.917, 2023, 2023.083, 2023.167,
    2023.25, 2023.333, 2023.417, 2023.5, 2023.583, 2023.667, 2023.75, 2023.833,
    2023.917, 2024 ;
}
