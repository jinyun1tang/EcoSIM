netcdf Lake_grid_20230221 {
dimensions:
	ncol = 1 ;
	nrow = 1 ;
	ngrid = 1 ;
	ntopou = 1 ;
	nlevs = 20 ;
variables:
	float ALATG(ngrid) ;
		ALATG:long_name = "Latitude" ;
		ALATG:units = "degrees north" ;
	float ALTIG(ngrid) ;
		ALTIG:long_name = "Altitude above sea-level" ;
		ALTIG:units = "m" ;
	float ATCAG(ngrid) ;
		ATCAG:long_name = "Mean annual temperaure" ;
		ATCAG:units = "oC" ;
	byte IDTBLG(ngrid) ;
		IDTBLG:long_name = "Water table flag" ;
		IDTBLG:units = "none" ;
		IDTBLG:flags = "0=No water table,1=Natural stationary water table,2=Natural mobile water table,3=Artificial stationary water table,4=Artificial mobile water table" ;
	float OXYEG(ngrid) ;
		OXYEG:long_name = "Atmospheric O2" ;
		OXYEG:units = "ppm" ;
	float Z2GEG(ngrid) ;
		Z2GEG:long_name = "Atmospheric N2" ;
		Z2GEG:units = "ppm" ;
	float CO2EIG(ngrid) ;
		CO2EIG:long_name = "Atmospheric CO2" ;
		CO2EIG:units = "ppm" ;
	float CH4EG(ngrid) ;
		CH4EG:long_name = "Atmospheric CH4" ;
		CH4EG:units = "ppm" ;
	float Z2OEG(ngrid) ;
		Z2OEG:long_name = "Atmospheric N2O" ;
		Z2OEG:units = "ppm" ;
	float ZNH3EG(ngrid) ;
		ZNH3EG:long_name = "Atmospheric NH3" ;
		ZNH3EG:units = "ppm" ;
	byte IETYPG(ngrid) ;
		IETYPG:long_name = "Koppen climate zone" ;
		IETYPG:units = "none" ;
	byte IERSNG(ngrid) ;
		IERSNG:long_name = "Flag for erosion model" ;
		IERSNG:units = "none" ;
		IERSNG:flags = "-1=no change in elevation,0=freeze-thaw to change elevation,1=freeze-thaw plus erosion to change elevation,2=freeze-thaw plus SOC accumulation to change elevation,3=freeze-thaw plus SOC accumulation, plus erosion to change elevation" ;
	byte NCNG(ngrid) ;
		NCNG:long_name = "Flag for lateral connections between grid cells" ;
		NCNG:units = "none" ;
		NCNG:flags = "0=No lateral connnection,1=Along the west-east direction,2=Along the north-south direction,3=3D lateral connection" ;
	float DTBLIG(ngrid) ;
		DTBLIG:long_name = "Depth of natural water table" ;
		DTBLIG:units = "m" ;
	float DTBLDIG(ngrid) ;
		DTBLDIG:long_name = "Depth of artificial water table" ;
		DTBLDIG:units = "m" ;
	float DTBLGG(ngrid) ;
		DTBLGG:long_name = "Slope of natural water table relative to landscape surface" ;
		DTBLGG:units = "none" ;
	float RCHQNG(ngrid) ;
		RCHQNG:long_name = "Boundary condition for North surface runoff" ;
		RCHQNG:units = "none" ;
		RCHQNG:flags = "varying between 0 and 1" ;
	float RCHQEG(ngrid) ;
		RCHQEG:long_name = "Boundary condition for East surface runoff" ;
		RCHQEG:units = "none" ;
		RCHQEG:flags = "varying between 0 and 1" ;
	float RCHQSG(ngrid) ;
		RCHQSG:long_name = "Boundary condition for S surface runoff" ;
		RCHQSG:units = "none" ;
		RCHQSG:flags = "varying between 0 and 1" ;
	float RCHQWG(ngrid) ;
		RCHQWG:long_name = "Boundary condition for W surface runoff" ;
		RCHQWG:units = "none" ;
		RCHQWG:flags = "varying between 0 and 1" ;
	float RCHGNUG(ngrid) ;
		RCHGNUG:long_name = "Bound condition for N subsurf flow" ;
		RCHGNUG:units = "none" ;
	float RCHGEUG(ngrid) ;
		RCHGEUG:long_name = "Bound condition for E subsurf flow" ;
		RCHGEUG:units = "none" ;
	float RCHGSUG(ngrid) ;
		RCHGSUG:long_name = "Bound condition for S subsurf flow" ;
		RCHGSUG:units = "none" ;
	float RCHGWUG(ngrid) ;
		RCHGWUG:long_name = "Bound condition for W subsurf flow" ;
		RCHGWUG:units = "none" ;
	float RCHGNTG(ngrid) ;
		RCHGNTG:long_name = "North edge distance to water table" ;
		RCHGNTG:units = "m" ;
	float RCHGETG(ngrid) ;
		RCHGETG:long_name = "East edge distance to water table" ;
		RCHGETG:units = "m" ;
	float RCHGSTG(ngrid) ;
		RCHGSTG:long_name = "South edge distance to water table" ;
		RCHGSTG:units = "m" ;
	float RCHGWTG(ngrid) ;
		RCHGWTG:long_name = "West edge distance to water table" ;
		RCHGWTG:units = "m" ;
	float RCHGDG(ngrid) ;
		RCHGDG:long_name = "Lower boundary conditions for water flow" ;
		RCHGDG:units = "none" ;
		RCHGDG:flags = "varying between 0 and 1" ;
	float DHI(ngrid, ncol) ;
	float DVI(ngrid, nrow) ;
	int topo_grid(ntopou) ;
		topo_grid:long_name = "grid ID of the topo unit" ;
		topo_grid:units = "none" ;
	byte NH1(ntopou) ;
		NH1:long_name = "Starting column from the west" ;
		NH1:units = "none" ;
	byte NH2(ntopou) ;
		NH2:long_name = "Ending column at the east" ;
		NH2:units = "none" ;
	byte NV1(ntopou) ;
		NV1:long_name = "Starting row from the north" ;
		NV1:units = "none" ;
	byte NV2(ntopou) ;
		NV2:long_name = "Ending row at the south" ;
		NV2:units = "none" ;
	float ASPX(ntopou) ;
		ASPX:long_name = "Aspect" ;
		ASPX:units = "degrees" ;
	float SL0(ntopou) ;
		SL0:long_name = "Slope" ;
		SL0:units = "degrees" ;
	float DPTHSX(ntopou) ;
		DPTHSX:long_name = "Initial snowpack depth" ;
		DPTHSX:units = "m" ;
	float PSIFC(ntopou) ;
		PSIFC:long_name = "Water potential at field capacity" ;
		PSIFC:units = "MPa" ;
	float PSIWP(ntopou) ;
		PSIWP:long_name = "Water potential at wilting point" ;
		PSIWP:units = "MPa" ;
	float ALBS(ntopou) ;
		ALBS:long_name = "Wet soil albedo" ;
		ALBS:units = "none" ;
	float PH0(ntopou) ;
		PH0:long_name = "Litter pH" ;
		PH0:units = "none" ;
	float RSCf(ntopou) ;
		RSCf:long_name = "C in surface fine litter" ;
		RSCf:units = "gC m-2" ;
	float RSNf(ntopou) ;
		RSNf:long_name = "N in surface fine litter" ;
		RSNf:units = "gN m-2" ;
	float RSPf(ntopou) ;
		RSPf:long_name = "P in surface fine litter" ;
		RSPf:units = "gP m-2" ;
	float RSCw(ntopou) ;
		RSCw:long_name = "C in surface woody litter" ;
		RSCw:units = "gC m-2" ;
	float RSNw(ntopou) ;
		RSNw:long_name = "N in surface woody litter" ;
		RSNw:units = "gN m-2" ;
	float RSPw(ntopou) ;
		RSPw:long_name = "P in surface woody litter" ;
		RSPw:units = "gP m-2" ;
	float RSCm(ntopou) ;
		RSCm:long_name = "C in manure" ;
		RSCm:units = "gC m-2" ;
	float RSNm(ntopou) ;
		RSNm:long_name = "N in manure" ;
		RSNm:units = "gN m-2" ;
	float RSPm(ntopou) ;
		RSPm:long_name = "P in manure" ;
		RSPm:units = "gP m-2" ;
	byte IXTYP1(ntopou) ;
		IXTYP1:long_name = "plant surface fine litter type" ;
		IXTYP1:units = "none" ;
		IXTYP1:flags = "1=maize,2=wheat,3=soybean,4=new straw,5=old straw,6=compost,7=green manure,8=new deciduos forest,9=new coniferous forest,10=old deciduous forest,11=old coniferous forest,12=default" ;
	byte IXTYP2(ntopou) ;
		IXTYP2:long_name = "manure surface litter type" ;
		IXTYP2:units = "none" ;
		IXTYP2:flags = "1=ruminant,2=non ruminant,3=others" ;
	byte NUI(ntopou) ;
		NUI:long_name = "Initial layer number of soil surface layer" ;
		NUI:units = "none" ;
		NUI:flags = "usually is 1" ;
	byte NJ(ntopou) ;
		NJ:long_name = "Layer number of maximum rooting layer" ;
		NJ:units = "none" ;
	byte NL1(ntopou) ;
		NL1:long_name = "Number of additional layers below NJ with data in file" ;
		NL1:units = "none" ;
	byte NL2(ntopou) ;
		NL2:long_name = "Number of additional layers below NJ without data in file" ;
		NL2:units = "none" ;
	byte ISOILR(ntopou) ;
		ISOILR:long_name = "Flag for soil profile type" ;
		ISOILR:units = "none" ;
		ISOILR:flags = "0=natural,1=reconstructed" ;
	float CDPTH(ntopou, nlevs) ;
		CDPTH:FillValue = -999.9 ;
		CDPTH:long_name = "Depth to bottom of soil layer" ;
		CDPTH:units = "m" ;
	float BKDSI(ntopou, nlevs) ;
		BKDSI:FillValue = -999.9 ;
		BKDSI:long_name = "Initial bulk density" ;
		BKDSI:units = "Mg m-3" ;
		BKDSI:flags = "0 for water" ;
	float FC(ntopou, nlevs) ;
		FC:FillValue = -999.9 ;
		FC:long_name = "Field capacity" ;
		FC:units = "m3 m-3" ;
	float WP(ntopou, nlevs) ;
		WP:FillValue = -999.9 ;
		WP:long_name = "Wilting point" ;
		WP:units = "m3 m-3" ;
	float SCNV(ntopou, nlevs) ;
		SCNV:FillValue = -999.9 ;
		SCNV:long_name = "Vertical hydraulic conductivity Ksat" ;
		SCNV:units = "mm h-1" ;
	float SCNH(ntopou, nlevs) ;
		SCNH:FillValue = -999.9 ;
		SCNH:long_name = "Lateral hydraulic conductivity Ksat" ;
		SCNH:units = "mm h-1" ;
	float CSAND(ntopou, nlevs) ;
		CSAND:FillValue = -999.9 ;
		CSAND:long_name = "Sand content" ;
		CSAND:units = "kg Mg-1" ;
	float CSILT(ntopou, nlevs) ;
		CSILT:FillValue = -999.9 ;
		CSILT:long_name = "Silt content" ;
		CSILT:units = "kg Mg-1" ;
	float FHOL(ntopou, nlevs) ;
		FHOL:FillValue = -999.9 ;
		FHOL:long_name = "Macropore fraction in the non-rock fraction of soil" ;
		FHOL:units = "none" ;
		FHOL:flags = "0-1" ;
	float ROCK(ntopou, nlevs) ;
		ROCK:FillValue = -999.9 ;
		ROCK:long_name = "Rock fraction of the whole soil" ;
		ROCK:units = "none" ;
		ROCK:flags = "0-1" ;
	float PH(ntopou, nlevs) ;
		PH:FillValue = -999.9 ;
		PH:long_name = "depth-resolved pH" ;
		PH:units = "none" ;
	float CEC(ntopou, nlevs) ;
		CEC:FillValue = -999.9 ;
		CEC:long_name = "Cation exchange capacity" ;
		CEC:units = "cmol kg soil-1" ;
	float AEC(ntopou, nlevs) ;
		AEC:FillValue = -999.9 ;
		AEC:long_name = "Anion exchange capacity" ;
		AEC:units = "cmol kg soil-1" ;
	float CORGC(ntopou, nlevs) ;
		CORGC:FillValue = -999.9 ;
		CORGC:long_name = "Total soil organic carbon" ;
		CORGC:units = "kg C/Mg soil" ;
	float CORGR(ntopou, nlevs) ;
		CORGR:FillValue = -999.9 ;
		CORGR:long_name = "POC (part of SOC)" ;
		CORGR:units = "kg C/Mg soil" ;
	float CORGN(ntopou, nlevs) ;
		CORGN:FillValue = -999.9 ;
		CORGN:long_name = "Total soil organic nitrogen" ;
		CORGN:units = "g N/Mg soil" ;
	float CORGP(ntopou, nlevs) ;
		CORGP:FillValue = -999.9 ;
		CORGP:long_name = "Total soil organic phosphorus" ;
		CORGP:units = "g P/Mg soil" ;
	float CNH4(ntopou, nlevs) ;
		CNH4:FillValue = -999.9 ;
		CNH4:long_name = "Total soil NH4 concentration" ;
		CNH4:units = "gN/Mg soil" ;
	float CNO3(ntopou, nlevs) ;
		CNO3:FillValue = -999.9 ;
		CNO3:long_name = "Total soil NO3 concentration" ;
		CNO3:units = "gN/Mg soil" ;
	float CPO4(ntopou, nlevs) ;
		CPO4:FillValue = -999.9 ;
		CPO4:long_name = "Total soil H2PO4 concentration" ;
		CPO4:units = "gP/Mg soil" ;
	float CAL(ntopou, nlevs) ;
		CAL:FillValue = -999.9 ;
		CAL:long_name = "Soluble soil Al content" ;
		CAL:units = "g Al/Mg soil" ;
	float CFE(ntopou, nlevs) ;
		CFE:FillValue = -999.9 ;
		CFE:long_name = "Soluble soil Fe content" ;
		CFE:units = "g Fe/Mg soil" ;
	float CCA(ntopou, nlevs) ;
		CCA:FillValue = -999.9 ;
		CCA:long_name = "Soluble soil Ca content" ;
		CCA:units = "g Ca/Mg soil" ;
	float CMG(ntopou, nlevs) ;
		CMG:FillValue = -999.9 ;
		CMG:long_name = "Soluble soil MG content" ;
		CMG:units = "g MG/Mg soil" ;
	float CNA(ntopou, nlevs) ;
		CNA:FillValue = -999.9 ;
		CNA:long_name = "Soluble soil Na content" ;
		CNA:units = "g Na/Mg soil" ;
	float CKA(ntopou, nlevs) ;
		CKA:FillValue = -999.9 ;
		CKA:long_name = "Soluble soil K content" ;
		CKA:units = "g K/Mg soil" ;
	float CSO4(ntopou, nlevs) ;
		CSO4:FillValue = -999.9 ;
		CSO4:long_name = "Soluble soil SO4 content" ;
		CSO4:units = "g S/Mg soil" ;
	float CCL(ntopou, nlevs) ;
		CCL:FillValue = -999.9 ;
		CCL:long_name = "Soluble soil Cl content" ;
		CCL:units = "g Cl/Mg soil" ;
	float CALPO(ntopou, nlevs) ;
		CALPO:FillValue = -999.9 ;
		CALPO:long_name = "Soil AlPO4 content" ;
		CALPO:units = "g P/Mg soil" ;
	float CFEPO(ntopou, nlevs) ;
		CFEPO:FillValue = -999.9 ;
		CFEPO:long_name = "Soil FePO4 content" ;
		CFEPO:units = "g P/Mg soil" ;
	float CCAPD(ntopou, nlevs) ;
		CCAPD:FillValue = -999.9 ;
		CCAPD:long_name = "Soil CaHPO4 content" ;
		CCAPD:units = "g P/Mg soil" ;
	float CCAPH(ntopou, nlevs) ;
		CCAPH:FillValue = -999.9 ;
		CCAPH:long_name = "Soil apatite content" ;
		CCAPH:units = "g P/Mg soil" ;
	float CALOH(ntopou, nlevs) ;
		CALOH:FillValue = -999.9 ;
		CALOH:long_name = "Soil Al(OH)3 content" ;
		CALOH:units = "g Al/Mg soil" ;
	float CFEOH(ntopou, nlevs) ;
		CFEOH:FillValue = -999.9 ;
		CFEOH:long_name = "Soil Fe(OH)3 content" ;
		CFEOH:units = "g Fe/Mg soil" ;
	float CCACO(ntopou, nlevs) ;
		CCACO:FillValue = -999.9 ;
		CCACO:long_name = "Soil CaCO3 content" ;
		CCACO:units = "g Ca/Mg soil" ;
	float CCASO(ntopou, nlevs) ;
		CCASO:FillValue = -999.9 ;
		CCASO:long_name = "Soil CaSO4 content" ;
		CCASO:units = "g Ca/Mg soil" ;
	float GKC4(ntopou, nlevs) ;
		GKC4:FillValue = -999.9 ;
		GKC4:long_name = "Ca-NH4 Gapon selectivity coefficient" ;
		GKC4:units = "none" ;
	float GKCH(ntopou, nlevs) ;
		GKCH:FillValue = -999.9 ;
		GKCH:long_name = "Ca-H Gapon selectivity coefficient" ;
		GKCH:units = "none" ;
	float GKCA(ntopou, nlevs) ;
		GKCA:FillValue = -999.9 ;
		GKCA:long_name = "Ca-Al Gapon selectivity coefficient" ;
		GKCA:units = "none" ;
	float GKCM(ntopou, nlevs) ;
		GKCM:FillValue = -999.9 ;
		GKCM:long_name = "Ca-Mg Gapon selectivity coefficient" ;
		GKCM:units = "none" ;
	float GKCN(ntopou, nlevs) ;
		GKCN:FillValue = -999.9 ;
		GKCN:long_name = "Ca-Na Gapon selectivity coefficient" ;
		GKCN:units = "none" ;
	float GKCK(ntopou, nlevs) ;
		GKCK:FillValue = -999.9 ;
		GKCK:long_name = "Ca-K Gapon selectivity coefficient" ;
		GKCK:units = "none" ;
	float THW(ntopou, nlevs) ;
		THW:FillValue = -999.9 ;
		THW:long_name = "Initial soil water content" ;
		THW:units = "m3/m3" ;
	float THI(ntopou, nlevs) ;
		THI:FillValue = -999.9 ;
		THI:long_name = "Initial soil ice content" ;
		THI:units = "m3/m3" ;
	float RSCfL(ntopou, nlevs) ;
		RSCfL:FillValue = -999.9 ;
		RSCfL:long_name = "Initial fine litter C" ;
		RSCfL:units = "gC m-2" ;
	float RSNfL(ntopou, nlevs) ;
		RSNfL:FillValue = -999.9 ;
		RSNfL:long_name = "Initial fine litter N" ;
		RSNfL:units = "gN m-2" ;
	float RSPfL(ntopou, nlevs) ;
		RSPfL:FillValue = -999.9 ;
		RSPfL:long_name = "Initial fine litter P" ;
		RSPfL:units = "gP m-2" ;
	float RSCwL(ntopou, nlevs) ;
		RSCwL:FillValue = -999.9 ;
		RSCwL:long_name = "Initial woody litter C" ;
		RSCwL:units = "gC m-2" ;
	float RSNwL(ntopou, nlevs) ;
		RSNwL:FillValue = -999.9 ;
		RSNwL:long_name = "Initial woody litter N" ;
		RSNwL:units = "gN m-2" ;
	float RSPwL(ntopou, nlevs) ;
		RSPwL:FillValue = -999.9 ;
		RSPwL:long_name = "Initial woody litter P" ;
		RSPwL:units = "gP m-2" ;
	float RSCmL(ntopou, nlevs) ;
		RSCmL:FillValue = -999.9 ;
		RSCmL:long_name = "Initial manure liter C" ;
		RSCmL:units = "gC m-2" ;
	float RSNmL(ntopou, nlevs) ;
		RSNmL:FillValue = -999.9 ;
		RSNmL:long_name = "Initial manure litter N" ;
		RSNmL:units = "gN m-2" ;
	float RSPmL(ntopou, nlevs) ;
		RSPmL:FillValue = -999.9 ;
		RSPmL:long_name = "Initial manure litter P" ;
		RSPmL:units = "gP m-2" ;
	int NHW ;
	int NHE ;
	int NVN ;
	int NVS ;

// global attributes:
		:description = "Grid input data created on 2023/02/21/18:26:08" ;
data:

 ALATG = 69.1 ;

 ALTIG = 130 ;

 ATCAG = -8 ;

 IDTBLG = 1 ;

 OXYEG = 210000 ;

 Z2GEG = 780000 ;

 CO2EIG = 326 ;

 CH4EG = 1.8 ;

 Z2OEG = 0.3 ;

 ZNH3EG = 0.005 ;

 IETYPG = 62 ;

 IERSNG = 0 ;

 NCNG = 1 ;

 DTBLIG = 3 ;

 DTBLDIG = 100 ;

 DTBLGG = 0 ;

 RCHQNG = 0 ;

 RCHQEG = 0 ;

 RCHQSG = 0 ;

 RCHQWG = 0 ;

 RCHGNUG = 0 ;

 RCHGEUG = 0 ;

 RCHGSUG = 0 ;

 RCHGWUG = 0 ;

 RCHGNTG = 0 ;

 RCHGETG = 0 ;

 RCHGSTG = 0 ;

 RCHGWTG = 0 ;

 RCHGDG = 0 ;

 DHI =
  1 ;

 DVI =
  1 ;

 topo_grid = 1 ;

 NH1 = 1 ;

 NH2 = 1 ;

 NV1 = 1 ;

 NV2 = 1 ;

 ASPX = 90 ;

 SL0 = 1 ;

 DPTHSX = 0 ;

 PSIFC = -0.03 ;

 PSIWP = -1.5 ;

 ALBS = 0.12 ;

 PH0 = 3.72 ;

 RSCf = 0. ;

 RSNf = 0. ;

 RSPf = 0. ;

 RSCw = 0 ;

 RSNw = 0 ;

 RSPw = 0 ;

 RSCm = 0 ;

 RSNm = 0 ;

 RSPm = 0 ;

 IXTYP1 = 10 ;

 IXTYP2 = 0 ;

 NUI = 1 ;

 NJ = 16 ;

 NL1 = 0 ;

 NL2 = 0 ;

 ISOILR = 1 ;

 CDPTH =
  0.01, 0.05, 0.15, 0.3, 0.5, 0.7, 1.16, 1.52, 1.82, 2.12, 2.42, 2.72, 3.1, 3.5, 3.9, 4.3, -999, -999, 
    -999, -999 ;

 BKDSI =
  0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0,0.0,0.0,1.47,1.47, 1.47, 1.47, 1.47,1.47,
    1.47,1.47,1.47, -999 ;

 FC =
  -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -999 ;

 WP =
  -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -999 ;

 SCNV =
  -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -999 ;

 SCNH =
  -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -999 ;

 CSAND =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 319.71, 319.71, 319.71, 319.71, 330.14, 330.14, 330.14, 330.14, 180, -999 ;

 CSILT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 545.39, 545.39, 545.39, 545.39, 184.49, 184.49, 184.49, 184.49, 20,  -999 ;

 FHOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -999 ;

 ROCK =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -999 ;

 PH =
  6.0, 6.0, 6.0, 6.0, 5.77, 5.77, 5.77, 5.77, 5.8, 5.8, 5.8, 5.8, 4.35, 4.35, 4.35, 4.35, 4.35, 
    4.35, 4.35,  -999 ;

 CEC =
  5.8, 5.8, 5.8, 5.8, 5.77, 5.77, 5.77, 5.77, 5.8, 5.8, 5.8, 5.8, 4.35, 4.35, 4.35, 4.35, 4.35, 
    4.35, 4.35,  -999 ;

 AEC =
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3,  -999 ;

 CORGC =
   0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.6, 2.6, 2, 2, 2, 2, 3, 0.5, 0.5, -999 ;

 CORGR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -999 ;

 CORGN =
  -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -999 ;

 CORGP =
  -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -999 ;

 CNH4 =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 3, 1, 1, 1, 0, 0, 0, -999 ;

 CNO3 =
   0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 12, 12, 1, 1, 1, 0, 0, 0, -999 ;

 CPO4 =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 10, 10, 10, 10, 10, 10, 10, 10,  -999 ;

 CAL =
  -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -999 ;

 CFE =
  -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 0, 0, 0, 0, 0, 0, 0, 0, -999 ;

 CCA =
  40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 
    -999 ;

 CMG =
  0, 0, 0, 18, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -999 ;

 CNA =
  0, 0, 0, 0, 0, 0, 0, 0,0, 0, 0.07, 0.05, 0.05, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01,  -999 ;

 CKA =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -999 ;

 CSO4 =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 48, 48, 48, 48, 48, 48, 48, 48,  -999 ;

 CCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 35, 35, 35, 35, 35, 35, 35, 35,  -999 ;

 CALPO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 50, 50, 50, 50, 50, 50, 50, 50, -999 ;

 CFEPO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 50, 50, 50, 50, 50, 50, 50, 50,  -999 ;

 CCAPD =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -999 ;

 CCAPH =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -999 ;

 CALOH =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, -999 ;

 CFEOH =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000,  -999 ;

 CCACO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -999 ;

 CCASO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -999 ;

 GKC4 =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, -999 ;

 GKCH =
  0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25, -999 ;

 GKCA =
  0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25, -999 ;

 GKCM =
  0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 
    0.6, -999 ;

 GKCN =
  0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, -999 ;

 GKCK =
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, -999 ;

 THW =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, -999 ;

 THI =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -999 ;

 RSCfL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 60, 75, 75, 60, 60, 45, 45, 15, -999 ;

 RSNfL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.5, 2, 2.5, 2.5, 2, 2, 1.5, 1.5, 0.5,  -999 ;

 RSPfL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.15, 0.2, 0.25, 0.25, 0.2, 0.2, 0.15, 0.15, 0.05,  -999 ;

 RSCwL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -999 ;

 RSNwL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -999 ;

 RSPwL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -999 ;

 RSCmL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -999 ;

 RSNmL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -999 ;

 RSPmL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -999 ;

 NHW = 1 ;

 NHE = 1 ;

 NVN = 1 ;

 NVS = 1 ;
}
