netcdf RiceUSTWT_soilmgmt_20251017 {
dimensions:
	ntopou = 1 ;
	nchar1 = 10 ;
	nchart = 24 ;
	nfert = 12 ;
	nfire = 12 ;
	nirri = 24 ;
	nchari = 128 ;
	ncharf = 128 ;
	year = UNLIMITED ; // (9 currently)
	ntill = 367 ;
variables:
	int year(year) ;
		year:long_name = "year AD" ;
	int NH1(ntopou) ;
		NH1:long_name = "Starting column from the west for a topo unit" ;
		NH1:units = "None" ;
	int NV1(ntopou) ;
		NV1:long_name = "Ending column at the east for a topo unit" ;
		NV1:units = "None" ;
	int NH2(ntopou) ;
		NH2:long_name = "Starting row from the north  for a topo unit" ;
		NH2:units = "None" ;
	int NV2(ntopou) ;
		NV2:long_name = "Ending row at the south  for a topo unit" ;
		NV2:units = "None" ;
	char fertf(year, ntopou, nchar1) ;
		fertf:long_name = "Fertilization info for a topo unit" ;
	char tillf(year, ntopou, nchar1) ;
		tillf:long_name = "Tillage info for a topo unit" ;
	char irrigf(year, ntopou, nchar1) ;
		irrigf:long_name = "Irrigation info for a topo unit" ;
	char me2008t(ntill, nchart) ;
		me2008t:long_name = "Tillage file" ;
	char me2008f(nfert, ncharf) ;
		me2008f:long_name = "Fertilization file" ;
	char me2009t(ntill, nchart) ;
		me2009t:long_name = "Tillage file" ;
	char me2009f(nfert, ncharf) ;
		me2009f:long_name = "Fertilization file" ;
	char me2010t(ntill, nchart) ;
		me2010t:long_name = "Tillage file" ;
	char me2010f(nfert, ncharf) ;
		me2010f:long_name = "Fertilization file" ;
	char me2011t(ntill, nchart) ;
		me2011t:long_name = "Tillage file" ;
	char me2011f(nfert, ncharf) ;
		me2011f:long_name = "Fertilization file" ;
	char me2012t(ntill, nchart) ;
		me2012t:long_name = "Tillage file" ;
	char me2012f(nfert, ncharf) ;
		me2012f:long_name = "Fertilization file" ;
	char me2013t(ntill, nchart) ;
		me2013t:long_name = "Tillage file" ;
	char me2013f(nfert, ncharf) ;
		me2013f:long_name = "Fertilization file" ;
	char me2014t(ntill, nchart) ;
		me2014t:long_name = "Tillage file" ;
	char me2014f(nfert, ncharf) ;
		me2014f:long_name = "Fertilization file" ;
	char me2015t(ntill, nchart) ;
		me2015t:long_name = "Tillage file" ;
	char me2015f(nfert, ncharf) ;
		me2015f:long_name = "Fertilization file" ;
	char me2016t(ntill, nchart) ;
		me2016t:long_name = "Tillage file" ;
	char me2016f(nfert, ncharf) ;
		me2016f:long_name = "Fertilization file" ;

// global attributes:
		:description = "soil managment data created on 2025/10/17/14:17:38" ;
data:

 year = 2008, 2009, 2010, 2011, 2012, 2013, 2014, 2015, 2016 ;

 NH1 = 1 ;

 NV1 = 1 ;

 NH2 = 1 ;

 NV2 = 1 ;

 fertf =
  "me2008f   ",
  "me2009f   ",
  "me2010f   ",
  "me2011f   ",
  "me2012f   ",
  "me2013f   ",
  "me2014f   ",
  "me2015f   ",
  "me2016f   " ;

 tillf =
  "me2008t   ",
  "me2009t   ",
  "me2010t   ",
  "me2011t   ",
  "me2012t   ",
  "me2013t   ",
  "me2014t   ",
  "me2015t   ",
  "me2016t   " ;

 irrigf =
  "NO        ",
  "NO        ",
  "NO        ",
  "NO        ",
  "NO        ",
  "NO        ",
  "NO        ",
  "NO        ",
  "NO        " ;

 me2008t =
  "15042008,3,0.100000     ",
  "01012008,23,-0.038109   ",
  "02012008,23,-0.034537   ",
  "03012008,23,-0.022564   ",
  "04012008,23,-0.013089   ",
  "05012008,23,-0.000118   ",
  "06012008,23,0.016454    ",
  "07012008,23,0.032126    ",
  "08012008,23,0.048490    ",
  "09012008,23,0.063872    ",
  "10012008,23,0.075422    ",
  "11012008,23,0.078677    ",
  "12012008,23,0.059362    ",
  "13012008,23,-0.008862   ",
  "14012008,23,-0.011899   ",
  "15012008,23,-0.004444   ",
  "16012008,23,0.003782    ",
  "17012008,23,0.012654    ",
  "18012008,23,0.009703    ",
  "19012008,23,0.005267    ",
  "20012008,23,-0.008881   ",
  "21012008,23,-0.037573   ",
  "22012008,23,-0.050234   ",
  "23012008,23,-0.043063   ",
  "24012008,23,-0.041937   ",
  "25012008,23,-0.037378   ",
  "26012008,23,-0.047049   ",
  "27012008,23,-0.038154   ",
  "28012008,23,-0.022005   ",
  "29012008,23,-0.010380   ",
  "30012008,23,0.001907    ",
  "31012008,23,0.023682    ",
  "01022008,23,0.049754    ",
  "02022008,23,0.070001    ",
  "03022008,23,0.090982    ",
  "04022008,23,0.103071    ",
  "05022008,23,0.087203    ",
  "06022008,23,0.091535    ",
  "07022008,23,0.126270    ",
  "08022008,23,0.163879    ",
  "09022008,23,0.163995    ",
  "10022008,23,0.213966    ",
  "11022008,23,0.261250    ",
  "12022008,23,0.299344    ",
  "13022008,23,0.330978    ",
  "14022008,23,0.364927    ",
  "15022008,23,0.397005    ",
  "16022008,23,0.430211    ",
  "17022008,23,0.455278    ",
  "18022008,23,0.467270    ",
  "19022008,23,0.484453    ",
  "20022008,23,0.508662    ",
  "21022008,23,0.517489    ",
  "22022008,23,0.488402    ",
  "23022008,23,0.457380    ",
  "24022008,23,0.292324    ",
  "25022008,23,0.363061    ",
  "26022008,23,0.361424    ",
  "27022008,23,0.320250    ",
  "28022008,23,0.397981    ",
  "01032008,23,0.458944    ",
  "02032008,23,0.418215    ",
  "03032008,23,0.269184    ",
  "04032008,23,0.246186    ",
  "05032008,23,0.286214    ",
  "06032008,23,0.316155    ",
  "07032008,23,0.371833    ",
  "08032008,23,0.454486    ",
  "09032008,23,0.510722    ",
  "10032008,23,0.529212    ",
  "11032008,23,0.396981    ",
  "12032008,23,0.423723    ",
  "13032008,23,0.500635    ",
  "14032008,23,0.475087    ",
  "15032008,23,0.475213    ",
  "16032008,23,0.457957    ",
  "17032008,23,0.481331    ",
  "18032008,23,0.466208    ",
  "19032008,23,0.463040    ",
  "20032008,23,0.437906    ",
  "21032008,23,0.441005    ",
  "22032008,23,0.469302    ",
  "23032008,23,0.524950    ",
  "24032008,23,0.436865    ",
  "25032008,23,0.389392    ",
  "26032008,23,0.435268    ",
  "27032008,23,0.506161    ",
  "28032008,23,0.493184    ",
  "29032008,23,0.533187    ",
  "30032008,23,0.508249    ",
  "31032008,23,0.502213    ",
  "01042008,23,0.488758    ",
  "02042008,23,0.577268    ",
  "03042008,23,0.592769    ",
  "04042008,23,0.615710    ",
  "05042008,23,0.614634    ",
  "06042008,23,0.612474    ",
  "07042008,23,0.634504    ",
  "08042008,23,0.644609    ",
  "09042008,23,0.621917    ",
  "10042008,23,0.635469    ",
  "11042008,23,0.634212    ",
  "12042008,23,0.635348    ",
  "13042008,23,0.636040    ",
  "14042008,23,0.645279    ",
  "15042008,23,0.648161    ",
  "16042008,23,0.627282    ",
  "17042008,23,0.627654    ",
  "18042008,23,0.633149    ",
  "19042008,23,0.646116    ",
  "20042008,23,0.640339    ",
  "21042008,23,0.648886    ",
  "22042008,23,0.653484    ",
  "23042008,23,0.610469    ",
  "24042008,23,0.632584    ",
  "25042008,23,0.643199    ",
  "26042008,23,0.652221    ",
  "27042008,23,0.658123    ",
  "28042008,23,0.668196    ",
  "29042008,23,0.676573    ",
  "30042008,23,0.683138    ",
  "01052008,23,0.686051    ",
  "02052008,23,0.695184    ",
  "03052008,23,0.704566    ",
  "04052008,23,0.706750    ",
  "05052008,23,0.709785    ",
  "06052008,23,0.717195    ",
  "07052008,23,0.720420    ",
  "08052008,23,0.723999    ",
  "09052008,23,0.728789    ",
  "10052008,23,0.731310    ",
  "11052008,23,0.732646    ",
  "12052008,23,0.725639    ",
  "13052008,23,0.720732    ",
  "14052008,23,0.724953    ",
  "15052008,23,0.730385    ",
  "16052008,23,0.731917    ",
  "17052008,23,0.737256    ",
  "18052008,23,0.743844    ",
  "19052008,23,0.751158    ",
  "20052008,23,0.758095    ",
  "21052008,23,0.764110    ",
  "22052008,23,0.772042    ",
  "23052008,23,0.774328    ",
  "24052008,23,0.783056    ",
  "25052008,23,0.785966    ",
  "26052008,23,0.778862    ",
  "27052008,23,0.777089    ",
  "28052008,23,0.768920    ",
  "29052008,23,0.771525    ",
  "30052008,23,0.785805    ",
  "31052008,23,0.802054    ",
  "01062008,23,0.816616    ",
  "02062008,23,0.830151    ",
  "03062008,23,0.841173    ",
  "04062008,23,0.851095    ",
  "05062008,23,0.861676    ",
  "06062008,23,0.873647    ",
  "07062008,23,0.883889    ",
  "08062008,23,0.893863    ",
  "09062008,23,0.905796    ",
  "10062008,23,0.914991    ",
  "11062008,23,0.923106    ",
  "12062008,23,0.806238    ",
  "13062008,23,0.589215    ",
  "14062008,23,0.101968    ",
  "15062008,23,-0.047320   ",
  "16062008,23,-0.053493   ",
  "17062008,23,-0.058756   ",
  "18062008,23,-0.057460   ",
  "19062008,23,-0.054845   ",
  "20062008,23,-0.061472   ",
  "21062008,23,-0.061128   ",
  "22062008,23,-0.056406   ",
  "23062008,23,-0.058857   ",
  "24062008,23,-0.044052   ",
  "25062008,23,-0.034997   ",
  "26062008,23,-0.032462   ",
  "27062008,23,-0.040039   ",
  "28062008,23,-0.044495   ",
  "29062008,23,-0.039912   ",
  "30062008,23,-0.034943   ",
  "01072008,23,-0.033777   ",
  "02072008,23,-0.032675   ",
  "03072008,23,-0.025429   ",
  "04072008,23,-0.019372   ",
  "05072008,23,-0.018008   ",
  "06072008,23,-0.015563   ",
  "07072008,23,-0.013608   ",
  "08072008,23,-0.028238   ",
  "09072008,23,-0.024172   ",
  "10072008,23,-0.018614   ",
  "11072008,23,-0.012971   ",
  "12072008,23,-0.003401   ",
  "13072008,23,0.002416    ",
  "14072008,23,0.000637    ",
  "15072008,23,-0.002413   ",
  "16072008,23,0.004379    ",
  "17072008,23,0.011109    ",
  "18072008,23,-0.003409   ",
  "19072008,23,-0.016766   ",
  "20072008,23,-0.031040   ",
  "21072008,23,-0.046582   ",
  "22072008,23,-0.070196   ",
  "23072008,23,-0.081960   ",
  "24072008,23,-0.146491   ",
  "25072008,23,-0.142168   ",
  "26072008,23,-0.138946   ",
  "27072008,23,-0.135727   ",
  "28072008,23,-0.132527   ",
  "29072008,23,-0.135403   ",
  "30072008,23,-0.137387   ",
  "31072008,23,-0.136588   ",
  "01082008,23,-0.136146   ",
  "02082008,23,-0.136016   ",
  "03082008,23,-0.135949   ",
  "04082008,23,-0.133109   ",
  "05082008,23,-0.130990   ",
  "06082008,23,-0.119439   ",
  "07082008,23,-0.123665   ",
  "08082008,23,-0.105511   ",
  "09082008,23,-0.101767   ",
  "10082008,23,-0.120952   ",
  "11082008,23,-0.109214   ",
  "12082008,23,-0.097563   ",
  "13082008,23,-0.095074   ",
  "14082008,23,-0.091981   ",
  "15082008,23,-0.094910   ",
  "16082008,23,-0.095380   ",
  "17082008,23,-0.093442   ",
  "18082008,23,-0.090215   ",
  "19082008,23,-0.086568   ",
  "20082008,23,-0.080672   ",
  "21082008,23,-0.080641   ",
  "22082008,23,-0.079274   ",
  "23082008,23,-0.077559   ",
  "24082008,23,-0.075271   ",
  "25082008,23,-0.074742   ",
  "26082008,23,-0.074262   ",
  "27082008,23,-0.072627   ",
  "28082008,23,-0.071035   ",
  "29082008,23,-0.067350   ",
  "30082008,23,-0.061547   ",
  "31082008,23,-0.059029   ",
  "01092008,23,-0.061018   ",
  "02092008,23,-0.062945   ",
  "03092008,23,-0.059135   ",
  "04092008,23,-0.055240   ",
  "05092008,23,-0.050484   ",
  "06092008,23,-0.044076   ",
  "07092008,23,-0.037188   ",
  "08092008,23,-0.034385   ",
  "09092008,23,-0.032871   ",
  "10092008,23,-0.037047   ",
  "11092008,23,-0.045285   ",
  "12092008,23,-0.055190   ",
  "13092008,23,-0.063886   ",
  "14092008,23,-0.080345   ",
  "15092008,23,-0.083851   ",
  "16092008,23,-0.073666   ",
  "17092008,23,-0.064057   ",
  "18092008,23,-0.049606   ",
  "19092008,23,-0.032421   ",
  "20092008,23,-0.012718   ",
  "21092008,23,0.011387    ",
  "22092008,23,0.032395    ",
  "23092008,23,0.088956    ",
  "24092008,23,0.192164    ",
  "25092008,23,0.319732    ",
  "26092008,23,0.416502    ",
  "27092008,23,0.468357    ",
  "28092008,23,0.535777    ",
  "29092008,23,0.593238    ",
  "30092008,23,0.633095    ",
  "01102008,23,0.664745    ",
  "02102008,23,0.672718    ",
  "03102008,23,0.702911    ",
  "04102008,23,0.729606    ",
  "05102008,23,0.748276    ",
  "06102008,23,0.688100    ",
  "07102008,23,0.682408    ",
  "08102008,23,0.693319    ",
  "09102008,23,0.706946    ",
  "10102008,23,0.714335    ",
  "11102008,23,0.723891    ",
  "12102008,23,0.608851    ",
  "13102008,23,0.653566    ",
  "14102008,23,0.479721    ",
  "15102008,23,0.446501    ",
  "16102008,23,0.500156    ",
  "17102008,23,0.427139    ",
  "18102008,23,0.471641    ",
  "19102008,23,0.621757    ",
  "20102008,23,0.503566    ",
  "21102008,23,0.611329    ",
  "22102008,23,0.571275    ",
  "23102008,23,0.543100    ",
  "24102008,23,0.503513    ",
  "25102008,23,0.550927    ",
  "26102008,23,0.514848    ",
  "27102008,23,0.547614    ",
  "28102008,23,0.491941    ",
  "29102008,23,0.396572    ",
  "30102008,23,0.374722    ",
  "31102008,23,0.294525    ",
  "01112008,23,0.217186    ",
  "02112008,23,0.151774    ",
  "03112008,23,0.128795    ",
  "04112008,23,0.103370    ",
  "05112008,23,0.069799    ",
  "06112008,23,0.184739    ",
  "07112008,23,0.200704    ",
  "08112008,23,0.165795    ",
  "09112008,23,0.129922    ",
  "10112008,23,0.064125    ",
  "11112008,23,0.053992    ",
  "12112008,23,0.046074    ",
  "13112008,23,0.164706    ",
  "14112008,23,0.133610    ",
  "15112008,23,0.101361    ",
  "16112008,23,0.124900    ",
  "17112008,23,0.069150    ",
  "18112008,23,0.049310    ",
  "19112008,23,0.005761    ",
  "20112008,23,0.386353    ",
  "21112008,23,0.155456    ",
  "22112008,23,0.015251    ",
  "23112008,23,-0.032184   ",
  "24112008,23,-0.068163   ",
  "25112008,23,-0.090485   ",
  "26112008,23,-0.087537   ",
  "27112008,23,-0.085009   ",
  "28112008,23,-0.102536   ",
  "29112008,23,-0.038977   ",
  "30112008,23,-0.020066   ",
  "01122008,23,-0.018299   ",
  "02122008,23,-0.033905   ",
  "03122008,23,-0.058786   ",
  "04122008,23,-0.078480   ",
  "05122008,23,-0.076164   ",
  "06122008,23,-0.074780   ",
  "07122008,23,-0.087493   ",
  "08122008,23,-0.071236   ",
  "09122008,23,-0.066845   ",
  "10122008,23,-0.067947   ",
  "11122008,23,-0.072111   ",
  "12122008,23,-0.071376   ",
  "13122008,23,-0.068235   ",
  "14122008,23,-0.068893   ",
  "15122008,23,-0.063309   ",
  "16122008,23,-0.065697   ",
  "17122008,23,-0.062278   ",
  "18122008,23,-0.061292   ",
  "19122008,23,-0.061507   ",
  "20122008,23,-0.063499   ",
  "21122008,23,-0.064303   ",
  "22122008,23,-0.075734   ",
  "23122008,23,-0.069499   ",
  "24122008,23,-0.057310   ",
  "25122008,23,-0.049512   ",
  "26122008,23,-0.041759   ",
  "27122008,23,-0.045208   ",
  "28122008,23,-0.047354   ",
  "29122008,23,-0.049188   ",
  "30122008,23,-0.047971   ",
  "31122008,23,-0.044181   ",
  "                        " ;

 me2008f =
  "16042008  0  0  0  0  5.82829  0  1.23291  0  0  0  0  0  0  0  0  0  0  0  0  0.02  0.76  0  0  1  0  0                        ",
  "07062008  0  0  0  0  0  0  5.04371  0  0  0  0  0  0  0  0  0  0  0  0  0.02  0.76  0  0  1  0  0                              ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                " ;

 me2009t =
  "15042009,3,0.100000     ",
  "01012009,23,-0.038109   ",
  "02012009,23,-0.034537   ",
  "03012009,23,-0.022564   ",
  "04012009,23,-0.013089   ",
  "05012009,23,-0.000118   ",
  "06012009,23,0.016454    ",
  "07012009,23,0.032126    ",
  "08012009,23,0.048490    ",
  "09012009,23,0.063872    ",
  "10012009,23,0.075422    ",
  "11012009,23,0.078677    ",
  "12012009,23,0.059362    ",
  "13012009,23,-0.008862   ",
  "14012009,23,-0.011899   ",
  "15012009,23,-0.004444   ",
  "16012009,23,0.003782    ",
  "17012009,23,0.012654    ",
  "18012009,23,0.009703    ",
  "19012009,23,0.005267    ",
  "20012009,23,-0.008881   ",
  "21012009,23,-0.037573   ",
  "22012009,23,-0.050234   ",
  "23012009,23,-0.043063   ",
  "24012009,23,-0.041937   ",
  "25012009,23,-0.037378   ",
  "26012009,23,-0.047049   ",
  "27012009,23,-0.038154   ",
  "28012009,23,-0.022005   ",
  "29012009,23,-0.010380   ",
  "30012009,23,0.001907    ",
  "31012009,23,0.023682    ",
  "01022009,23,0.049754    ",
  "02022009,23,0.070001    ",
  "03022009,23,0.090982    ",
  "04022009,23,0.103071    ",
  "05022009,23,0.087203    ",
  "06022009,23,0.091535    ",
  "07022009,23,0.126270    ",
  "08022009,23,0.163879    ",
  "09022009,23,0.163995    ",
  "10022009,23,0.213966    ",
  "11022009,23,0.261250    ",
  "12022009,23,0.299344    ",
  "13022009,23,0.330978    ",
  "14022009,23,0.364927    ",
  "15022009,23,0.397005    ",
  "16022009,23,0.430211    ",
  "17022009,23,0.455278    ",
  "18022009,23,0.467270    ",
  "19022009,23,0.484453    ",
  "20022009,23,0.508662    ",
  "21022009,23,0.517489    ",
  "22022009,23,0.488402    ",
  "23022009,23,0.457380    ",
  "24022009,23,0.292324    ",
  "25022009,23,0.363061    ",
  "26022009,23,0.361424    ",
  "27022009,23,0.320250    ",
  "28022009,23,0.397981    ",
  "01032009,23,0.458944    ",
  "02032009,23,0.418215    ",
  "03032009,23,0.269184    ",
  "04032009,23,0.246186    ",
  "05032009,23,0.286214    ",
  "06032009,23,0.316155    ",
  "07032009,23,0.371833    ",
  "08032009,23,0.454486    ",
  "09032009,23,0.510722    ",
  "10032009,23,0.529212    ",
  "11032009,23,0.396981    ",
  "12032009,23,0.423723    ",
  "13032009,23,0.500635    ",
  "14032009,23,0.475087    ",
  "15032009,23,0.475213    ",
  "16032009,23,0.457957    ",
  "17032009,23,0.481331    ",
  "18032009,23,0.466208    ",
  "19032009,23,0.463040    ",
  "20032009,23,0.437906    ",
  "21032009,23,0.441005    ",
  "22032009,23,0.469302    ",
  "23032009,23,0.524950    ",
  "24032009,23,0.436865    ",
  "25032009,23,0.389392    ",
  "26032009,23,0.435268    ",
  "27032009,23,0.506161    ",
  "28032009,23,0.493184    ",
  "29032009,23,0.533187    ",
  "30032009,23,0.508249    ",
  "31032009,23,0.502213    ",
  "01042009,23,0.488758    ",
  "02042009,23,0.577268    ",
  "03042009,23,0.592769    ",
  "04042009,23,0.615710    ",
  "05042009,23,0.614634    ",
  "06042009,23,0.612474    ",
  "07042009,23,0.634504    ",
  "08042009,23,0.644609    ",
  "09042009,23,0.621917    ",
  "10042009,23,0.635469    ",
  "11042009,23,0.634212    ",
  "12042009,23,0.635348    ",
  "13042009,23,0.636040    ",
  "14042009,23,0.645279    ",
  "15042009,23,0.648161    ",
  "16042009,23,0.627282    ",
  "17042009,23,0.627654    ",
  "18042009,23,0.633149    ",
  "19042009,23,0.646116    ",
  "20042009,23,0.640339    ",
  "21042009,23,0.648886    ",
  "22042009,23,0.653484    ",
  "23042009,23,0.610469    ",
  "24042009,23,0.632584    ",
  "25042009,23,0.643199    ",
  "26042009,23,0.652221    ",
  "27042009,23,0.658123    ",
  "28042009,23,0.668196    ",
  "29042009,23,0.676573    ",
  "30042009,23,0.683138    ",
  "01052009,23,0.686051    ",
  "02052009,23,0.695184    ",
  "03052009,23,0.704566    ",
  "04052009,23,0.706750    ",
  "05052009,23,0.709785    ",
  "06052009,23,0.717195    ",
  "07052009,23,0.720420    ",
  "08052009,23,0.723999    ",
  "09052009,23,0.728789    ",
  "10052009,23,0.731310    ",
  "11052009,23,0.732646    ",
  "12052009,23,0.725639    ",
  "13052009,23,0.720732    ",
  "14052009,23,0.724953    ",
  "15052009,23,0.730385    ",
  "16052009,23,0.731917    ",
  "17052009,23,0.737256    ",
  "18052009,23,0.743844    ",
  "19052009,23,0.751158    ",
  "20052009,23,0.758095    ",
  "21052009,23,0.764110    ",
  "22052009,23,0.772042    ",
  "23052009,23,0.774328    ",
  "24052009,23,0.783056    ",
  "25052009,23,0.785966    ",
  "26052009,23,0.778862    ",
  "27052009,23,0.777089    ",
  "28052009,23,0.768920    ",
  "29052009,23,0.771525    ",
  "30052009,23,0.785805    ",
  "31052009,23,0.802054    ",
  "01062009,23,0.816616    ",
  "02062009,23,0.830151    ",
  "03062009,23,0.841173    ",
  "04062009,23,0.851095    ",
  "05062009,23,0.861676    ",
  "06062009,23,0.873647    ",
  "07062009,23,0.883889    ",
  "08062009,23,0.893863    ",
  "09062009,23,0.905796    ",
  "10062009,23,0.914991    ",
  "11062009,23,0.923106    ",
  "12062009,23,0.806238    ",
  "13062009,23,0.589215    ",
  "14062009,23,0.101968    ",
  "15062009,23,-0.047320   ",
  "16062009,23,-0.053493   ",
  "17062009,23,-0.058756   ",
  "18062009,23,-0.057460   ",
  "19062009,23,-0.054845   ",
  "20062009,23,-0.061472   ",
  "21062009,23,-0.061128   ",
  "22062009,23,-0.056406   ",
  "23062009,23,-0.058857   ",
  "24062009,23,-0.044052   ",
  "25062009,23,-0.034997   ",
  "26062009,23,-0.032462   ",
  "27062009,23,-0.040039   ",
  "28062009,23,-0.044495   ",
  "29062009,23,-0.039912   ",
  "30062009,23,-0.034943   ",
  "01072009,23,-0.033777   ",
  "02072009,23,-0.032675   ",
  "03072009,23,-0.025429   ",
  "04072009,23,-0.019372   ",
  "05072009,23,-0.018008   ",
  "06072009,23,-0.015563   ",
  "07072009,23,-0.013608   ",
  "08072009,23,-0.028238   ",
  "09072009,23,-0.024172   ",
  "10072009,23,-0.018614   ",
  "11072009,23,-0.012971   ",
  "12072009,23,-0.003401   ",
  "13072009,23,0.002416    ",
  "14072009,23,0.000637    ",
  "15072009,23,-0.002413   ",
  "16072009,23,0.004379    ",
  "17072009,23,0.011109    ",
  "18072009,23,-0.003409   ",
  "19072009,23,-0.016766   ",
  "20072009,23,-0.031040   ",
  "21072009,23,-0.046582   ",
  "22072009,23,-0.070196   ",
  "23072009,23,-0.081960   ",
  "24072009,23,-0.146491   ",
  "25072009,23,-0.142168   ",
  "26072009,23,-0.138946   ",
  "27072009,23,-0.135727   ",
  "28072009,23,-0.132527   ",
  "29072009,23,-0.135403   ",
  "30072009,23,-0.137387   ",
  "31072009,23,-0.136588   ",
  "01082009,23,-0.136146   ",
  "02082009,23,-0.136016   ",
  "03082009,23,-0.135949   ",
  "04082009,23,-0.133109   ",
  "05082009,23,-0.130990   ",
  "06082009,23,-0.119439   ",
  "07082009,23,-0.123665   ",
  "08082009,23,-0.105511   ",
  "09082009,23,-0.101767   ",
  "10082009,23,-0.120952   ",
  "11082009,23,-0.109214   ",
  "12082009,23,-0.097563   ",
  "13082009,23,-0.095074   ",
  "14082009,23,-0.091981   ",
  "15082009,23,-0.094910   ",
  "16082009,23,-0.095380   ",
  "17082009,23,-0.093442   ",
  "18082009,23,-0.090215   ",
  "19082009,23,-0.086568   ",
  "20082009,23,-0.080672   ",
  "21082009,23,-0.080641   ",
  "22082009,23,-0.079274   ",
  "23082009,23,-0.077559   ",
  "24082009,23,-0.075271   ",
  "25082009,23,-0.074742   ",
  "26082009,23,-0.074262   ",
  "27082009,23,-0.072627   ",
  "28082009,23,-0.071035   ",
  "29082009,23,-0.067350   ",
  "30082009,23,-0.061547   ",
  "31082009,23,-0.059029   ",
  "01092009,23,-0.061018   ",
  "02092009,23,-0.062945   ",
  "03092009,23,-0.059135   ",
  "04092009,23,-0.055240   ",
  "05092009,23,-0.050484   ",
  "06092009,23,-0.044076   ",
  "07092009,23,-0.037188   ",
  "08092009,23,-0.034385   ",
  "09092009,23,-0.032871   ",
  "10092009,23,-0.037047   ",
  "11092009,23,-0.045285   ",
  "12092009,23,-0.055190   ",
  "13092009,23,-0.063886   ",
  "14092009,23,-0.080345   ",
  "15092009,23,-0.083851   ",
  "16092009,23,-0.073666   ",
  "17092009,23,-0.064057   ",
  "18092009,23,-0.049606   ",
  "19092009,23,-0.032421   ",
  "20092009,23,-0.012718   ",
  "21092009,23,0.011387    ",
  "22092009,23,0.032395    ",
  "23092009,23,0.088956    ",
  "24092009,23,0.192164    ",
  "25092009,23,0.319732    ",
  "26092009,23,0.416502    ",
  "27092009,23,0.468357    ",
  "28092009,23,0.535777    ",
  "29092009,23,0.593238    ",
  "30092009,23,0.633095    ",
  "01102009,23,0.664745    ",
  "02102009,23,0.672718    ",
  "03102009,23,0.702911    ",
  "04102009,23,0.729606    ",
  "05102009,23,0.748276    ",
  "06102009,23,0.688100    ",
  "07102009,23,0.682408    ",
  "08102009,23,0.693319    ",
  "09102009,23,0.706946    ",
  "10102009,23,0.714335    ",
  "11102009,23,0.723891    ",
  "12102009,23,0.608851    ",
  "13102009,23,0.653566    ",
  "14102009,23,0.479721    ",
  "15102009,23,0.446501    ",
  "16102009,23,0.500156    ",
  "17102009,23,0.427139    ",
  "18102009,23,0.471641    ",
  "19102009,23,0.621757    ",
  "20102009,23,0.503566    ",
  "21102009,23,0.611329    ",
  "22102009,23,0.571275    ",
  "23102009,23,0.543100    ",
  "24102009,23,0.503513    ",
  "25102009,23,0.550927    ",
  "26102009,23,0.514848    ",
  "27102009,23,0.547614    ",
  "28102009,23,0.491941    ",
  "29102009,23,0.396572    ",
  "30102009,23,0.374722    ",
  "31102009,23,0.294525    ",
  "01112009,23,0.217186    ",
  "02112009,23,0.151774    ",
  "03112009,23,0.128795    ",
  "04112009,23,0.103370    ",
  "05112009,23,0.069799    ",
  "06112009,23,0.184739    ",
  "07112009,23,0.200704    ",
  "08112009,23,0.165795    ",
  "09112009,23,0.129922    ",
  "10112009,23,0.064125    ",
  "11112009,23,0.053992    ",
  "12112009,23,0.046074    ",
  "13112009,23,0.164706    ",
  "14112009,23,0.133610    ",
  "15112009,23,0.101361    ",
  "16112009,23,0.124900    ",
  "17112009,23,0.069150    ",
  "18112009,23,0.049310    ",
  "19112009,23,0.005761    ",
  "20112009,23,0.386353    ",
  "21112009,23,0.155456    ",
  "22112009,23,0.015251    ",
  "23112009,23,-0.032184   ",
  "24112009,23,-0.068163   ",
  "25112009,23,-0.090485   ",
  "26112009,23,-0.087537   ",
  "27112009,23,-0.085009   ",
  "28112009,23,-0.102536   ",
  "29112009,23,-0.038977   ",
  "30112009,23,-0.020066   ",
  "01122009,23,-0.018299   ",
  "02122009,23,-0.033905   ",
  "03122009,23,-0.058786   ",
  "04122009,23,-0.078480   ",
  "05122009,23,-0.076164   ",
  "06122009,23,-0.074780   ",
  "07122009,23,-0.087493   ",
  "08122009,23,-0.071236   ",
  "09122009,23,-0.066845   ",
  "10122009,23,-0.067947   ",
  "11122009,23,-0.072111   ",
  "12122009,23,-0.071376   ",
  "13122009,23,-0.068235   ",
  "14122009,23,-0.068893   ",
  "15122009,23,-0.063309   ",
  "16122009,23,-0.065697   ",
  "17122009,23,-0.062278   ",
  "18122009,23,-0.061292   ",
  "19122009,23,-0.061507   ",
  "20122009,23,-0.063499   ",
  "21122009,23,-0.064303   ",
  "22122009,23,-0.075734   ",
  "23122009,23,-0.069499   ",
  "24122009,23,-0.057310   ",
  "25122009,23,-0.049512   ",
  "26122009,23,-0.041759   ",
  "27122009,23,-0.045208   ",
  "28122009,23,-0.047354   ",
  "29122009,23,-0.049188   ",
  "30122009,23,-0.047971   ",
  "31122009,23,-0.044181   ",
  "                        " ;

 me2009f =
  "16042009  0  0  0  0  5.82829  0  1.23291  0  0  0  0  0  0  0  0  0  0  0  0  0.02  0.76  0  0  1  0  0                        ",
  "07062009  0  0  0  0  0  0  5.04371  0  0  0  0  0  0  0  0  0  0  0  0  0.02  0.76  0  0  1  0  0                              ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                " ;

 me2010t =
  "15042010,3,0.100000     ",
  "01012010,23,-0.038109   ",
  "02012010,23,-0.034537   ",
  "03012010,23,-0.022564   ",
  "04012010,23,-0.013089   ",
  "05012010,23,-0.000118   ",
  "06012010,23,0.016454    ",
  "07012010,23,0.032126    ",
  "08012010,23,0.048490    ",
  "09012010,23,0.063872    ",
  "10012010,23,0.075422    ",
  "11012010,23,0.078677    ",
  "12012010,23,0.059362    ",
  "13012010,23,-0.008862   ",
  "14012010,23,-0.011899   ",
  "15012010,23,-0.004444   ",
  "16012010,23,0.003782    ",
  "17012010,23,0.012654    ",
  "18012010,23,0.009703    ",
  "19012010,23,0.005267    ",
  "20012010,23,-0.008881   ",
  "21012010,23,-0.037573   ",
  "22012010,23,-0.050234   ",
  "23012010,23,-0.043063   ",
  "24012010,23,-0.041937   ",
  "25012010,23,-0.037378   ",
  "26012010,23,-0.047049   ",
  "27012010,23,-0.038154   ",
  "28012010,23,-0.022005   ",
  "29012010,23,-0.010380   ",
  "30012010,23,0.001907    ",
  "31012010,23,0.023682    ",
  "01022010,23,0.049754    ",
  "02022010,23,0.070001    ",
  "03022010,23,0.090982    ",
  "04022010,23,0.103071    ",
  "05022010,23,0.087203    ",
  "06022010,23,0.091535    ",
  "07022010,23,0.126270    ",
  "08022010,23,0.163879    ",
  "09022010,23,0.163995    ",
  "10022010,23,0.213966    ",
  "11022010,23,0.261250    ",
  "12022010,23,0.299344    ",
  "13022010,23,0.330978    ",
  "14022010,23,0.364927    ",
  "15022010,23,0.397005    ",
  "16022010,23,0.430211    ",
  "17022010,23,0.455278    ",
  "18022010,23,0.467270    ",
  "19022010,23,0.484453    ",
  "20022010,23,0.508662    ",
  "21022010,23,0.517489    ",
  "22022010,23,0.488402    ",
  "23022010,23,0.457380    ",
  "24022010,23,0.292324    ",
  "25022010,23,0.363061    ",
  "26022010,23,0.361424    ",
  "27022010,23,0.320250    ",
  "28022010,23,0.397981    ",
  "01032010,23,0.458944    ",
  "02032010,23,0.418215    ",
  "03032010,23,0.269184    ",
  "04032010,23,0.246186    ",
  "05032010,23,0.286214    ",
  "06032010,23,0.316155    ",
  "07032010,23,0.371833    ",
  "08032010,23,0.454486    ",
  "09032010,23,0.510722    ",
  "10032010,23,0.529212    ",
  "11032010,23,0.396981    ",
  "12032010,23,0.423723    ",
  "13032010,23,0.500635    ",
  "14032010,23,0.475087    ",
  "15032010,23,0.475213    ",
  "16032010,23,0.457957    ",
  "17032010,23,0.481331    ",
  "18032010,23,0.466208    ",
  "19032010,23,0.463040    ",
  "20032010,23,0.437906    ",
  "21032010,23,0.441005    ",
  "22032010,23,0.469302    ",
  "23032010,23,0.524950    ",
  "24032010,23,0.436865    ",
  "25032010,23,0.389392    ",
  "26032010,23,0.435268    ",
  "27032010,23,0.506161    ",
  "28032010,23,0.493184    ",
  "29032010,23,0.533187    ",
  "30032010,23,0.508249    ",
  "31032010,23,0.502213    ",
  "01042010,23,0.488758    ",
  "02042010,23,0.577268    ",
  "03042010,23,0.592769    ",
  "04042010,23,0.615710    ",
  "05042010,23,0.614634    ",
  "06042010,23,0.612474    ",
  "07042010,23,0.634504    ",
  "08042010,23,0.644609    ",
  "09042010,23,0.621917    ",
  "10042010,23,0.635469    ",
  "11042010,23,0.634212    ",
  "12042010,23,0.635348    ",
  "13042010,23,0.636040    ",
  "14042010,23,0.645279    ",
  "15042010,23,0.648161    ",
  "16042010,23,0.627282    ",
  "17042010,23,0.627654    ",
  "18042010,23,0.633149    ",
  "19042010,23,0.646116    ",
  "20042010,23,0.640339    ",
  "21042010,23,0.648886    ",
  "22042010,23,0.653484    ",
  "23042010,23,0.610469    ",
  "24042010,23,0.632584    ",
  "25042010,23,0.643199    ",
  "26042010,23,0.652221    ",
  "27042010,23,0.658123    ",
  "28042010,23,0.668196    ",
  "29042010,23,0.676573    ",
  "30042010,23,0.683138    ",
  "01052010,23,0.686051    ",
  "02052010,23,0.695184    ",
  "03052010,23,0.704566    ",
  "04052010,23,0.706750    ",
  "05052010,23,0.709785    ",
  "06052010,23,0.717195    ",
  "07052010,23,0.720420    ",
  "08052010,23,0.723999    ",
  "09052010,23,0.728789    ",
  "10052010,23,0.731310    ",
  "11052010,23,0.732646    ",
  "12052010,23,0.725639    ",
  "13052010,23,0.720732    ",
  "14052010,23,0.724953    ",
  "15052010,23,0.730385    ",
  "16052010,23,0.731917    ",
  "17052010,23,0.737256    ",
  "18052010,23,0.743844    ",
  "19052010,23,0.751158    ",
  "20052010,23,0.758095    ",
  "21052010,23,0.764110    ",
  "22052010,23,0.772042    ",
  "23052010,23,0.774328    ",
  "24052010,23,0.783056    ",
  "25052010,23,0.785966    ",
  "26052010,23,0.778862    ",
  "27052010,23,0.777089    ",
  "28052010,23,0.768920    ",
  "29052010,23,0.771525    ",
  "30052010,23,0.785805    ",
  "31052010,23,0.802054    ",
  "01062010,23,0.816616    ",
  "02062010,23,0.830151    ",
  "03062010,23,0.841173    ",
  "04062010,23,0.851095    ",
  "05062010,23,0.861676    ",
  "06062010,23,0.873647    ",
  "07062010,23,0.883889    ",
  "08062010,23,0.893863    ",
  "09062010,23,0.905796    ",
  "10062010,23,0.914991    ",
  "11062010,23,0.923106    ",
  "12062010,23,0.806238    ",
  "13062010,23,0.589215    ",
  "14062010,23,0.101968    ",
  "15062010,23,-0.047320   ",
  "16062010,23,-0.053493   ",
  "17062010,23,-0.058756   ",
  "18062010,23,-0.057460   ",
  "19062010,23,-0.054845   ",
  "20062010,23,-0.061472   ",
  "21062010,23,-0.061128   ",
  "22062010,23,-0.056406   ",
  "23062010,23,-0.058857   ",
  "24062010,23,-0.044052   ",
  "25062010,23,-0.034997   ",
  "26062010,23,-0.032462   ",
  "27062010,23,-0.040039   ",
  "28062010,23,-0.044495   ",
  "29062010,23,-0.039912   ",
  "30062010,23,-0.034943   ",
  "01072010,23,-0.033777   ",
  "02072010,23,-0.032675   ",
  "03072010,23,-0.025429   ",
  "04072010,23,-0.019372   ",
  "05072010,23,-0.018008   ",
  "06072010,23,-0.015563   ",
  "07072010,23,-0.013608   ",
  "08072010,23,-0.028238   ",
  "09072010,23,-0.024172   ",
  "10072010,23,-0.018614   ",
  "11072010,23,-0.012971   ",
  "12072010,23,-0.003401   ",
  "13072010,23,0.002416    ",
  "14072010,23,0.000637    ",
  "15072010,23,-0.002413   ",
  "16072010,23,0.004379    ",
  "17072010,23,0.011109    ",
  "18072010,23,-0.003409   ",
  "19072010,23,-0.016766   ",
  "20072010,23,-0.031040   ",
  "21072010,23,-0.046582   ",
  "22072010,23,-0.070196   ",
  "23072010,23,-0.081960   ",
  "24072010,23,-0.092505   ",
  "25072010,23,-0.107267   ",
  "26072010,23,-0.099198   ",
  "27072010,23,-0.090727   ",
  "28072010,23,-0.133817   ",
  "29072010,23,-0.185575   ",
  "30072010,23,-0.195236   ",
  "31072010,23,-0.198564   ",
  "01082010,23,-0.204108   ",
  "02082010,23,-0.208920   ",
  "03082010,23,-0.210394   ",
  "04082010,23,-0.209849   ",
  "05082010,23,-0.199309   ",
  "06082010,23,-0.195179   ",
  "07082010,23,-0.194606   ",
  "08082010,23,-0.191280   ",
  "09082010,23,-0.184636   ",
  "10082010,23,-0.173988   ",
  "11082010,23,-0.159428   ",
  "12082010,23,-0.157927   ",
  "13082010,23,-0.158758   ",
  "14082010,23,-0.159591   ",
  "15082010,23,-0.162515   ",
  "16082010,23,-0.165987   ",
  "17082010,23,-0.173605   ",
  "18082010,23,-0.178176   ",
  "19082010,23,-0.179925   ",
  "20082010,23,-0.180138   ",
  "21082010,23,-0.177886   ",
  "22082010,23,-0.177643   ",
  "23082010,23,-0.179066   ",
  "24082010,23,-0.179826   ",
  "25082010,23,-0.180197   ",
  "26082010,23,-0.177316   ",
  "27082010,23,-0.175894   ",
  "28082010,23,-0.174127   ",
  "29082010,23,-0.174212   ",
  "30082010,23,-0.173107   ",
  "31082010,23,-0.172571   ",
  "01092010,23,-0.169716   ",
  "02092010,23,-0.164402   ",
  "03092010,23,-0.156901   ",
  "04092010,23,-0.147774   ",
  "05092010,23,-0.135429   ",
  "06092010,23,-0.119235   ",
  "07092010,23,-0.098152   ",
  "08092010,23,-0.081738   ",
  "09092010,23,-0.068862   ",
  "10092010,23,-0.066122   ",
  "11092010,23,-0.061662   ",
  "12092010,23,-0.059523   ",
  "13092010,23,-0.061255   ",
  "14092010,23,-0.070973   ",
  "15092010,23,-0.101516   ",
  "16092010,23,-0.126684   ",
  "17092010,23,-0.144928   ",
  "18092010,23,-0.152865   ",
  "19092010,23,-0.155429   ",
  "20092010,23,-0.145150   ",
  "21092010,23,-0.101463   ",
  "22092010,23,-0.063937   ",
  "23092010,23,-0.031777   ",
  "24092010,23,0.004190    ",
  "25092010,23,0.025403    ",
  "26092010,23,0.050293    ",
  "27092010,23,0.104418    ",
  "28092010,23,0.180382    ",
  "29092010,23,0.252384    ",
  "30092010,23,0.336364    ",
  "01102010,23,0.410474    ",
  "02102010,23,0.459949    ",
  "03102010,23,0.507054    ",
  "04102010,23,0.539730    ",
  "05102010,23,0.567449    ",
  "06102010,23,0.594575    ",
  "07102010,23,0.618299    ",
  "08102010,23,0.634261    ",
  "09102010,23,0.648424    ",
  "10102010,23,0.658557    ",
  "11102010,23,0.669345    ",
  "12102010,23,0.688057    ",
  "13102010,23,0.701433    ",
  "14102010,23,0.711992    ",
  "15102010,23,0.720565    ",
  "16102010,23,0.732856    ",
  "17102010,23,0.745794    ",
  "18102010,23,0.747025    ",
  "19102010,23,0.749978    ",
  "20102010,23,0.756645    ",
  "21102010,23,0.765701    ",
  "22102010,23,0.771919    ",
  "23102010,23,0.774870    ",
  "24102010,23,0.749078    ",
  "25102010,23,0.699798    ",
  "26102010,23,0.694581    ",
  "27102010,23,0.730526    ",
  "28102010,23,0.727906    ",
  "29102010,23,0.727493    ",
  "30102010,23,0.738151    ",
  "31102010,23,0.703483    ",
  "01112010,23,0.712645    ",
  "02112010,23,0.701454    ",
  "03112010,23,0.709311    ",
  "04112010,23,0.715301    ",
  "05112010,23,0.733654    ",
  "06112010,23,0.724414    ",
  "07112010,23,0.602299    ",
  "08112010,23,0.287473    ",
  "09112010,23,0.021659    ",
  "10112010,23,-0.114912   ",
  "11112010,23,0.148253    ",
  "12112010,23,0.127369    ",
  "13112010,23,0.023126    ",
  "14112010,23,-0.096454   ",
  "15112010,23,-0.120652   ",
  "16112010,23,-0.119653   ",
  "17112010,23,-0.118340   ",
  "18112010,23,-0.115133   ",
  "19112010,23,-0.115804   ",
  "20112010,23,-0.112690   ",
  "21112010,23,-0.128144   ",
  "22112010,23,-0.114688   ",
  "23112010,23,-0.117478   ",
  "24112010,23,-0.103499   ",
  "25112010,23,-0.090653   ",
  "26112010,23,-0.093497   ",
  "27112010,23,-0.100647   ",
  "28112010,23,-0.102684   ",
  "29112010,23,-0.104441   ",
  "30112010,23,-0.120061   ",
  "01122010,23,-0.130599   ",
  "02122010,23,-0.136632   ",
  "03122010,23,-0.128023   ",
  "04122010,23,-0.117416   ",
  "05122010,23,-0.112534   ",
  "06122010,23,-0.112386   ",
  "07122010,23,-0.106286   ",
  "08122010,23,-0.103977   ",
  "09122010,23,-0.103498   ",
  "10122010,23,-0.097612   ",
  "11122010,23,-0.092653   ",
  "12122010,23,-0.090173   ",
  "13122010,23,-0.090024   ",
  "14122010,23,-0.093128   ",
  "15122010,23,-0.096371   ",
  "16122010,23,-0.094369   ",
  "17122010,23,-0.092407   ",
  "18122010,23,-0.089805   ",
  "19122010,23,-0.114012   ",
  "20122010,23,-0.113051   ",
  "21122010,23,-0.103441   ",
  "22122010,23,-0.100584   ",
  "23122010,23,-0.098421   ",
  "24122010,23,-0.101866   ",
  "25122010,23,-0.110460   ",
  "26122010,23,-0.108508   ",
  "27122010,23,-0.110615   ",
  "28122010,23,-0.109305   ",
  "29122010,23,-0.136172   ",
  "30122010,23,-0.108638   ",
  "31122010,23,-0.096857   ",
  "                        " ;

 me2010f =
  "16042010  0  0  0  0  5.82829  0  1.23291  0  0  0  0  0  0  0  0  0  0  0  0  0.02  0.76  0  0  1  0  0                        ",
  "07062010  0  0  0  0  0  0  5.04371  0  0  0  0  0  0  0  0  0  0  0  0  0.02  0.76  0  0  1  0  0                              ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                " ;

 me2011t =
  "22042011,3,0.100000     ",
  "01012011,23,-0.094235   ",
  "02012011,23,-0.107830   ",
  "03012011,23,-0.109069   ",
  "04012011,23,-0.106347   ",
  "05012011,23,-0.105509   ",
  "06012011,23,-0.104134   ",
  "07012011,23,-0.103435   ",
  "08012011,23,-0.099024   ",
  "09012011,23,-0.095117   ",
  "10012011,23,-0.091502   ",
  "11012011,23,-0.090494   ",
  "12012011,23,-0.090329   ",
  "13012011,23,-0.089773   ",
  "14012011,23,-0.090474   ",
  "15012011,23,-0.091043   ",
  "16012011,23,-0.092391   ",
  "17012011,23,-0.089260   ",
  "18012011,23,-0.090703   ",
  "19012011,23,-0.091411   ",
  "20012011,23,-0.084831   ",
  "21012011,23,-0.086301   ",
  "22012011,23,-0.085533   ",
  "23012011,23,-0.083232   ",
  "24012011,23,-0.085019   ",
  "25012011,23,-0.084419   ",
  "26012011,23,-0.081901   ",
  "27012011,23,-0.084951   ",
  "28012011,23,-0.085233   ",
  "29012011,23,-0.084367   ",
  "30012011,23,-0.089099   ",
  "31012011,23,-0.092800   ",
  "01022011,23,-0.091838   ",
  "02022011,23,-0.078000   ",
  "03022011,23,-0.079609   ",
  "04022011,23,-0.076587   ",
  "05022011,23,-0.077322   ",
  "06022011,23,-0.059411   ",
  "07022011,23,-0.046332   ",
  "08022011,23,-0.032999   ",
  "09022011,23,-0.000824   ",
  "10022011,23,0.003804    ",
  "11022011,23,0.012939    ",
  "12022011,23,0.020788    ",
  "13022011,23,0.021618    ",
  "14022011,23,0.027251    ",
  "15022011,23,0.025223    ",
  "16022011,23,0.016621    ",
  "17022011,23,0.015618    ",
  "18022011,23,0.008350    ",
  "19022011,23,0.005790    ",
  "20022011,23,0.030043    ",
  "21022011,23,0.030977    ",
  "22022011,23,0.040823    ",
  "23022011,23,0.038399    ",
  "24022011,23,0.038928    ",
  "25022011,23,0.019538    ",
  "26022011,23,0.029519    ",
  "27022011,23,0.038431    ",
  "28022011,23,0.042939    ",
  "01032011,23,0.043606    ",
  "02032011,23,0.039783    ",
  "03032011,23,0.045062    ",
  "04032011,23,0.048925    ",
  "05032011,23,0.049005    ",
  "06032011,23,0.025706    ",
  "07032011,23,0.033923    ",
  "08032011,23,0.046293    ",
  "09032011,23,0.043024    ",
  "10032011,23,0.039128    ",
  "11032011,23,0.039168    ",
  "12032011,23,0.047241    ",
  "13032011,23,0.057872    ",
  "14032011,23,0.060412    ",
  "15032011,23,0.047305    ",
  "16032011,23,0.038932    ",
  "17032011,23,0.071012    ",
  "18032011,23,0.055857    ",
  "19032011,23,0.025851    ",
  "20032011,23,0.019186    ",
  "21032011,23,0.038182    ",
  "22032011,23,0.050871    ",
  "23032011,23,0.035088    ",
  "24032011,23,0.026577    ",
  "25032011,23,0.027526    ",
  "26032011,23,0.024618    ",
  "27032011,23,0.030975    ",
  "28032011,23,0.038373    ",
  "29032011,23,0.046237    ",
  "30032011,23,0.055281    ",
  "31032011,23,0.064024    ",
  "01042011,23,0.070749    ",
  "02042011,23,0.099964    ",
  "03042011,23,0.166654    ",
  "04042011,23,0.201576    ",
  "05042011,23,0.240145    ",
  "06042011,23,0.289453    ",
  "07042011,23,0.307663    ",
  "08042011,23,0.332982    ",
  "09042011,23,0.385419    ",
  "10042011,23,0.442948    ",
  "11042011,23,0.332165    ",
  "12042011,23,0.356176    ",
  "13042011,23,0.359929    ",
  "14042011,23,0.393047    ",
  "15042011,23,0.377338    ",
  "16042011,23,0.388411    ",
  "17042011,23,0.423880    ",
  "18042011,23,0.442974    ",
  "19042011,23,0.506524    ",
  "20042011,23,0.553608    ",
  "21042011,23,0.554895    ",
  "22042011,23,0.586329    ",
  "23042011,23,0.599370    ",
  "24042011,23,0.596301    ",
  "25042011,23,0.612473    ",
  "26042011,23,0.608525    ",
  "27042011,23,0.592312    ",
  "28042011,23,0.600105    ",
  "29042011,23,0.615045    ",
  "30042011,23,0.615891    ",
  "01052011,23,0.625236    ",
  "02052011,23,0.637446    ",
  "03052011,23,0.595761    ",
  "04052011,23,0.579030    ",
  "05052011,23,0.584975    ",
  "06052011,23,0.588085    ",
  "07052011,23,0.611529    ",
  "08052011,23,0.616304    ",
  "09052011,23,0.626686    ",
  "10052011,23,0.633334    ",
  "11052011,23,0.640678    ",
  "12052011,23,0.194650    ",
  "13052011,23,-0.008509   ",
  "14052011,23,-0.031851   ",
  "15052011,23,-0.013144   ",
  "16052011,23,0.026067    ",
  "17052011,23,0.032322    ",
  "18052011,23,0.038552    ",
  "19052011,23,0.073222    ",
  "20052011,23,0.122975    ",
  "21052011,23,0.179024    ",
  "22052011,23,0.238112    ",
  "23052011,23,0.307918    ",
  "24052011,23,0.369668    ",
  "25052011,23,0.413362    ",
  "26052011,23,0.463987    ",
  "27052011,23,0.491772    ",
  "28052011,23,0.500629    ",
  "29052011,23,0.532076    ",
  "30052011,23,0.587699    ",
  "31052011,23,0.618948    ",
  "01062011,23,0.649912    ",
  "02062011,23,0.668850    ",
  "03062011,23,0.658900    ",
  "04062011,23,0.674964    ",
  "05062011,23,0.664921    ",
  "06062011,23,0.652154    ",
  "07062011,23,0.641688    ",
  "08062011,23,0.654160    ",
  "09062011,23,0.682994    ",
  "10062011,23,0.702901    ",
  "11062011,23,0.726304    ",
  "12062011,23,0.751641    ",
  "13062011,23,0.770815    ",
  "14062011,23,0.744899    ",
  "15062011,23,0.596871    ",
  "16062011,23,0.148627    ",
  "17062011,23,-0.015393   ",
  "18062011,23,-0.026939   ",
  "19062011,23,-0.035351   ",
  "20062011,23,-0.033742   ",
  "21062011,23,-0.016866   ",
  "22062011,23,-0.004805   ",
  "23062011,23,0.007931    ",
  "24062011,23,0.022666    ",
  "25062011,23,0.026453    ",
  "26062011,23,0.026097    ",
  "27062011,23,0.027457    ",
  "28062011,23,0.024072    ",
  "29062011,23,0.014732    ",
  "30062011,23,0.014923    ",
  "01072011,23,0.010109    ",
  "02072011,23,0.001850    ",
  "03072011,23,-0.009887   ",
  "04072011,23,-0.016085   ",
  "05072011,23,-0.022531   ",
  "06072011,23,-0.027144   ",
  "07072011,23,-0.028314   ",
  "08072011,23,-0.020040   ",
  "09072011,23,-0.073858   ",
  "10072011,23,-0.103802   ",
  "11072011,23,-0.128013   ",
  "12072011,23,-0.131239   ",
  "13072011,23,-0.131740   ",
  "14072011,23,-0.132747   ",
  "15072011,23,-0.129910   ",
  "16072011,23,-0.145424   ",
  "17072011,23,-0.127428   ",
  "18072011,23,-0.121208   ",
  "19072011,23,-0.117103   ",
  "20072011,23,-0.143456   ",
  "21072011,23,-0.150494   ",
  "22072011,23,-0.146644   ",
  "23072011,23,-0.107202   ",
  "24072011,23,-0.098202   ",
  "25072011,23,-0.091360   ",
  "26072011,23,-0.088904   ",
  "27072011,23,-0.085830   ",
  "28072011,23,-0.080586   ",
  "29072011,23,-0.074721   ",
  "30072011,23,-0.071551   ",
  "31072011,23,-0.075238   ",
  "01082011,23,-0.078758   ",
  "02082011,23,-0.084558   ",
  "03082011,23,-0.093171   ",
  "04082011,23,-0.099484   ",
  "05082011,23,-0.105853   ",
  "06082011,23,-0.112429   ",
  "07082011,23,-0.117541   ",
  "08082011,23,-0.122111   ",
  "09082011,23,-0.127418   ",
  "10082011,23,-0.132746   ",
  "11082011,23,-0.133897   ",
  "12082011,23,-0.135965   ",
  "13082011,23,-0.140234   ",
  "14082011,23,-0.140876   ",
  "15082011,23,-0.141472   ",
  "16082011,23,-0.143867   ",
  "17082011,23,-0.143481   ",
  "18082011,23,-0.141218   ",
  "19082011,23,-0.141598   ",
  "20082011,23,-0.141080   ",
  "21082011,23,-0.133035   ",
  "22082011,23,-0.128485   ",
  "23082011,23,-0.129128   ",
  "24082011,23,-0.129809   ",
  "25082011,23,-0.129375   ",
  "26082011,23,-0.130082   ",
  "27082011,23,-0.131088   ",
  "28082011,23,-0.131650   ",
  "29082011,23,-0.125343   ",
  "30082011,23,-0.112597   ",
  "31082011,23,-0.101377   ",
  "01092011,23,-0.088799   ",
  "02092011,23,-0.075527   ",
  "03092011,23,-0.062414   ",
  "04092011,23,-0.049647   ",
  "05092011,23,-0.036721   ",
  "06092011,23,-0.010582   ",
  "07092011,23,0.036619    ",
  "08092011,23,0.097133    ",
  "09092011,23,0.135046    ",
  "10092011,23,0.182451    ",
  "11092011,23,0.258942    ",
  "12092011,23,0.300848    ",
  "13092011,23,0.332834    ",
  "14092011,23,0.360257    ",
  "15092011,23,0.406300    ",
  "16092011,23,0.465074    ",
  "17092011,23,0.522081    ",
  "18092011,23,0.556124    ",
  "19092011,23,0.561490    ",
  "20092011,23,0.564229    ",
  "21092011,23,0.570980    ",
  "22092011,23,0.595659    ",
  "23092011,23,0.598457    ",
  "24092011,23,0.595642    ",
  "25092011,23,0.566714    ",
  "26092011,23,0.566386    ",
  "27092011,23,0.564249    ",
  "28092011,23,0.557455    ",
  "29092011,23,0.556613    ",
  "30092011,23,0.559543    ",
  "01102011,23,0.564357    ",
  "02102011,23,0.555525    ",
  "03102011,23,0.548495    ",
  "04102011,23,0.547605    ",
  "05102011,23,0.544939    ",
  "06102011,23,0.544090    ",
  "07102011,23,0.543938    ",
  "08102011,23,0.544834    ",
  "09102011,23,0.546352    ",
  "10102011,23,0.539174    ",
  "11102011,23,0.546391    ",
  "12102011,23,0.545760    ",
  "13102011,23,0.545131    ",
  "14102011,23,0.545429    ",
  "15102011,23,0.545832    ",
  "16102011,23,0.544298    ",
  "17102011,23,0.532311    ",
  "18102011,23,0.520453    ",
  "19102011,23,0.544831    ",
  "20102011,23,0.545035    ",
  "21102011,23,0.550394    ",
  "22102011,23,0.548723    ",
  "23102011,23,0.545776    ",
  "24102011,23,0.589384    ",
  "25102011,23,0.571383    ",
  "26102011,23,0.502049    ",
  "27102011,23,0.583902    ",
  "28102011,23,0.644980    ",
  "29102011,23,0.541042    ",
  "30102011,23,0.620050    ",
  "31102011,23,0.511023    ",
  "01112011,23,0.467494    ",
  "02112011,23,0.554273    ",
  "03112011,23,0.680397    ",
  "04112011,23,0.680742    ",
  "05112011,23,0.680713    ",
  "06112011,23,0.680745    ",
  "07112011,23,0.680643    ",
  "08112011,23,0.678170    ",
  "09112011,23,0.285328    ",
  "10112011,23,-0.129377   ",
  "11112011,23,-0.164570   ",
  "12112011,23,-0.187369   ",
  "13112011,23,-0.203985   ",
  "14112011,23,-0.181652   ",
  "15112011,23,-0.157493   ",
  "16112011,23,-0.153234   ",
  "17112011,23,-0.153253   ",
  "18112011,23,-0.143611   ",
  "19112011,23,-0.133404   ",
  "20112011,23,-0.133637   ",
  "21112011,23,-0.125638   ",
  "22112011,23,-0.116935   ",
  "23112011,23,-0.112000   ",
  "24112011,23,-0.107185   ",
  "25112011,23,-0.100386   ",
  "26112011,23,-0.092940   ",
  "27112011,23,-0.090043   ",
  "28112011,23,-0.090766   ",
  "29112011,23,-0.092457   ",
  "30112011,23,-0.093839   ",
  "01122011,23,-0.088252   ",
  "02122011,23,-0.081859   ",
  "03122011,23,-0.078874   ",
  "04122011,23,-0.075556   ",
  "05122011,23,-0.081827   ",
  "06122011,23,-0.095580   ",
  "07122011,23,-0.106745   ",
  "08122011,23,-0.111539   ",
  "09122011,23,-0.114770   ",
  "10122011,23,-0.117553   ",
  "11122011,23,-0.120318   ",
  "12122011,23,-0.121014   ",
  "13122011,23,-0.122272   ",
  "14122011,23,-0.120183   ",
  "15122011,23,-0.122665   ",
  "16122011,23,-0.122196   ",
  "17122011,23,-0.123278   ",
  "18122011,23,-0.125164   ",
  "19122011,23,-0.124179   ",
  "20122011,23,-0.124263   ",
  "21122011,23,-0.124768   ",
  "22122011,23,-0.111815   ",
  "23122011,23,-0.117160   ",
  "24122011,23,-0.118412   ",
  "25122011,23,-0.120258   ",
  "26122011,23,-0.122216   ",
  "27122011,23,-0.123074   ",
  "28122011,23,-0.120478   ",
  "29122011,23,-0.115227   ",
  "30122011,23,-0.109849   ",
  "31122011,23,-0.104020   ",
  "                        " ;

 me2011f =
  "22042011  0  0  0  0  5.82829  0  1.23291  0  0  0  0  0  0  0  0  0  0  0  0  0.02  0.76  0  0  1  0  0                        ",
  "14062011  0  0  0  0  0  0  6.72495  0  0  0  0  0  0  0  0  0  0  0  0  0.02  0.76  0  0  1  0  0                              ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                " ;

 me2012t =
  "17052012,3,0.100000     ",
  "01012012,23,-0.105201   ",
  "02012012,23,-0.106448   ",
  "03012012,23,-0.108551   ",
  "04012012,23,-0.111640   ",
  "05012012,23,-0.115970   ",
  "06012012,23,-0.119548   ",
  "07012012,23,-0.117728   ",
  "08012012,23,-0.113389   ",
  "09012012,23,-0.117701   ",
  "10012012,23,-0.120473   ",
  "11012012,23,-0.123072   ",
  "12012012,23,-0.125206   ",
  "13012012,23,-0.128139   ",
  "14012012,23,-0.130284   ",
  "15012012,23,-0.138061   ",
  "16012012,23,-0.120377   ",
  "17012012,23,-0.148355   ",
  "18012012,23,-0.149585   ",
  "19012012,23,-0.151498   ",
  "20012012,23,-0.153051   ",
  "21012012,23,-0.159215   ",
  "22012012,23,-0.139726   ",
  "23012012,23,-0.145382   ",
  "24012012,23,-0.142451   ",
  "25012012,23,-0.135820   ",
  "26012012,23,-0.126342   ",
  "27012012,23,-0.121452   ",
  "28012012,23,-0.129024   ",
  "29012012,23,-0.125551   ",
  "30012012,23,-0.125264   ",
  "31012012,23,-0.124969   ",
  "01022012,23,-0.119827   ",
  "02022012,23,-0.117299   ",
  "03022012,23,-0.115925   ",
  "04022012,23,-0.113387   ",
  "05022012,23,-0.111237   ",
  "06022012,23,-0.103229   ",
  "07022012,23,-0.100426   ",
  "08022012,23,-0.085513   ",
  "09022012,23,-0.068266   ",
  "10022012,23,-0.055352   ",
  "11022012,23,-0.048128   ",
  "12022012,23,-0.041800   ",
  "13022012,23,-0.042496   ",
  "14022012,23,-0.030402   ",
  "15022012,23,-0.023004   ",
  "16022012,23,-0.014571   ",
  "17022012,23,-0.009881   ",
  "18022012,23,-0.007157   ",
  "19022012,23,-0.002025   ",
  "20022012,23,0.002564    ",
  "21022012,23,0.006452    ",
  "22022012,23,0.009820    ",
  "23022012,23,0.023735    ",
  "24022012,23,0.080361    ",
  "25022012,23,0.120120    ",
  "26022012,23,0.116336    ",
  "27022012,23,0.142005    ",
  "28022012,23,0.206679    ",
  "29022012,23,0.156039    ",
  "01032012,23,0.126056    ",
  "02032012,23,0.176398    ",
  "03032012,23,0.207096    ",
  "04032012,23,0.210984    ",
  "05032012,23,0.222554    ",
  "06032012,23,0.254279    ",
  "07032012,23,0.315744    ",
  "08032012,23,0.360228    ",
  "09032012,23,0.366314    ",
  "10032012,23,0.351408    ",
  "11032012,23,0.378925    ",
  "12032012,23,0.393782    ",
  "13032012,23,0.358209    ",
  "14032012,23,0.077856    ",
  "15032012,23,0.009552    ",
  "16032012,23,0.013544    ",
  "17032012,23,-0.005192   ",
  "18032012,23,0.003708    ",
  "19032012,23,0.040979    ",
  "20032012,23,0.063577    ",
  "21032012,23,0.062020    ",
  "22032012,23,0.082809    ",
  "23032012,23,0.131483    ",
  "24032012,23,0.146308    ",
  "25032012,23,0.040432    ",
  "26032012,23,0.053915    ",
  "27032012,23,0.027738    ",
  "28032012,23,-0.002002   ",
  "29032012,23,0.008309    ",
  "30032012,23,0.013579    ",
  "31032012,23,0.017433    ",
  "01042012,23,0.052403    ",
  "02042012,23,0.058761    ",
  "03042012,23,0.089589    ",
  "04042012,23,0.147127    ",
  "05042012,23,0.183510    ",
  "06042012,23,0.216727    ",
  "07042012,23,0.230040    ",
  "08042012,23,0.133823    ",
  "09042012,23,0.138786    ",
  "10042012,23,0.096970    ",
  "11042012,23,0.126927    ",
  "12042012,23,0.152616    ",
  "13042012,23,0.147007    ",
  "14042012,23,0.152600    ",
  "15042012,23,0.119268    ",
  "16042012,23,0.120631    ",
  "17042012,23,0.120190    ",
  "18042012,23,0.136719    ",
  "19042012,23,0.158398    ",
  "20042012,23,0.166017    ",
  "21042012,23,0.180313    ",
  "22042012,23,0.183307    ",
  "23042012,23,0.120315    ",
  "24042012,23,0.072983    ",
  "25042012,23,0.070830    ",
  "26042012,23,0.084157    ",
  "27042012,23,0.117844    ",
  "28042012,23,0.013917    ",
  "29042012,23,0.018837    ",
  "30042012,23,0.109352    ",
  "01052012,23,-0.008568   ",
  "02052012,23,-0.001628   ",
  "03052012,23,-0.013411   ",
  "04052012,23,-0.034504   ",
  "05052012,23,-0.106638   ",
  "06052012,23,0.103369    ",
  "07052012,23,0.140520    ",
  "08052012,23,0.097718    ",
  "09052012,23,0.144962    ",
  "10052012,23,0.065868    ",
  "11052012,23,0.143387    ",
  "12052012,23,0.109310    ",
  "13052012,23,-0.043669   ",
  "14052012,23,-0.022794   ",
  "15052012,23,-0.095247   ",
  "16052012,23,-0.100925   ",
  "17052012,23,-0.110499   ",
  "18052012,23,-0.062222   ",
  "19052012,23,0.018660    ",
  "20052012,23,0.067242    ",
  "21052012,23,-0.068689   ",
  "22052012,23,-0.159169   ",
  "23052012,23,-0.126147   ",
  "24052012,23,-0.090294   ",
  "25052012,23,-0.056101   ",
  "26052012,23,-0.003171   ",
  "27052012,23,0.069545    ",
  "28052012,23,0.149690    ",
  "29052012,23,0.220433    ",
  "30052012,23,0.278967    ",
  "31052012,23,0.325274    ",
  "01062012,23,0.367209    ",
  "02062012,23,0.439316    ",
  "03062012,23,0.496366    ",
  "04062012,23,0.553331    ",
  "05062012,23,0.601096    ",
  "06062012,23,0.617691    ",
  "07062012,23,0.646141    ",
  "08062012,23,0.672477    ",
  "09062012,23,0.697878    ",
  "10062012,23,0.718934    ",
  "11062012,23,0.739201    ",
  "12062012,23,0.752350    ",
  "13062012,23,0.760814    ",
  "14062012,23,0.773788    ",
  "15062012,23,0.789435    ",
  "16062012,23,0.759104    ",
  "17062012,23,0.389899    ",
  "18062012,23,-0.058687   ",
  "19062012,23,-0.084999   ",
  "20062012,23,-0.094473   ",
  "21062012,23,-0.115012   ",
  "22062012,23,-0.105293   ",
  "23062012,23,-0.077255   ",
  "24062012,23,-0.056921   ",
  "25062012,23,-0.062310   ",
  "26062012,23,-0.059622   ",
  "27062012,23,-0.056520   ",
  "28062012,23,-0.059872   ",
  "29062012,23,-0.065075   ",
  "30062012,23,-0.065543   ",
  "01072012,23,-0.064871   ",
  "02072012,23,-0.121876   ",
  "03072012,23,-0.162048   ",
  "04072012,23,-0.174045   ",
  "05072012,23,-0.171461   ",
  "06072012,23,-0.170778   ",
  "07072012,23,-0.172060   ",
  "08072012,23,-0.170116   ",
  "09072012,23,-0.167151   ",
  "10072012,23,-0.165487   ",
  "11072012,23,-0.164924   ",
  "12072012,23,-0.160904   ",
  "13072012,23,-0.155357   ",
  "14072012,23,-0.150742   ",
  "15072012,23,-0.147936   ",
  "16072012,23,-0.140848   ",
  "17072012,23,-0.135677   ",
  "18072012,23,-0.140307   ",
  "19072012,23,-0.142099   ",
  "20072012,23,-0.145753   ",
  "21072012,23,-0.154289   ",
  "22072012,23,-0.164564   ",
  "23072012,23,-0.170794   ",
  "24072012,23,-0.178675   ",
  "25072012,23,-0.185505   ",
  "26072012,23,-0.188334   ",
  "27072012,23,-0.186505   ",
  "28072012,23,-0.187739   ",
  "29072012,23,-0.191601   ",
  "30072012,23,-0.193579   ",
  "31072012,23,-0.192538   ",
  "01082012,23,-0.193404   ",
  "02082012,23,-0.196120   ",
  "03082012,23,-0.195548   ",
  "04082012,23,-0.189319   ",
  "05082012,23,-0.189511   ",
  "06082012,23,-0.192003   ",
  "07082012,23,-0.193237   ",
  "08082012,23,-0.191143   ",
  "09082012,23,-0.192191   ",
  "10082012,23,-0.191521   ",
  "11082012,23,-0.186403   ",
  "12082012,23,-0.176984   ",
  "13082012,23,-0.173741   ",
  "14082012,23,-0.168879   ",
  "15082012,23,-0.163084   ",
  "16082012,23,-0.160549   ",
  "17082012,23,-0.158601   ",
  "18082012,23,-0.155569   ",
  "19082012,23,-0.154681   ",
  "20082012,23,-0.154213   ",
  "21082012,23,-0.153035   ",
  "22082012,23,-0.149330   ",
  "23082012,23,-0.146198   ",
  "24082012,23,-0.143233   ",
  "25082012,23,-0.141974   ",
  "26082012,23,-0.134882   ",
  "27082012,23,-0.138260   ",
  "28082012,23,-0.142406   ",
  "29082012,23,-0.146341   ",
  "30082012,23,-0.145564   ",
  "31082012,23,-0.141145   ",
  "01092012,23,-0.144015   ",
  "02092012,23,-0.148878   ",
  "03092012,23,-0.146523   ",
  "04092012,23,-0.142287   ",
  "05092012,23,-0.143223   ",
  "06092012,23,-0.141789   ",
  "07092012,23,-0.140240   ",
  "08092012,23,-0.137686   ",
  "09092012,23,-0.130858   ",
  "10092012,23,-0.129264   ",
  "11092012,23,-0.125908   ",
  "12092012,23,-0.126791   ",
  "13092012,23,-0.132907   ",
  "14092012,23,-0.135354   ",
  "15092012,23,-0.137461   ",
  "16092012,23,-0.138872   ",
  "17092012,23,-0.128912   ",
  "18092012,23,-0.115447   ",
  "19092012,23,-0.103349   ",
  "20092012,23,-0.092945   ",
  "21092012,23,-0.080034   ",
  "22092012,23,-0.067191   ",
  "23092012,23,-0.053054   ",
  "24092012,23,-0.026728   ",
  "25092012,23,0.017751    ",
  "26092012,23,0.073327    ",
  "27092012,23,0.128571    ",
  "28092012,23,0.183783    ",
  "29092012,23,0.239218    ",
  "30092012,23,0.271539    ",
  "01102012,23,0.294720    ",
  "02102012,23,0.318996    ",
  "03102012,23,0.360368    ",
  "04102012,23,0.417780    ",
  "05102012,23,0.451991    ",
  "06102012,23,0.470100    ",
  "07102012,23,0.499691    ",
  "08102012,23,0.540757    ",
  "09102012,23,0.565816    ",
  "10102012,23,0.586413    ",
  "11102012,23,0.617266    ",
  "12102012,23,0.661323    ",
  "13102012,23,0.680300    ",
  "14102012,23,0.684719    ",
  "15102012,23,0.690710    ",
  "16102012,23,0.703940    ",
  "17102012,23,0.724803    ",
  "18102012,23,0.749424    ",
  "19102012,23,0.764036    ",
  "20102012,23,0.770360    ",
  "21102012,23,0.788601    ",
  "22102012,23,0.789742    ",
  "23102012,23,0.766795    ",
  "24102012,23,0.759270    ",
  "25102012,23,0.771533    ",
  "26102012,23,0.764936    ",
  "27102012,23,0.756566    ",
  "28102012,23,0.760244    ",
  "29102012,23,0.763276    ",
  "30102012,23,0.762960    ",
  "31102012,23,0.767526    ",
  "01112012,23,0.773584    ",
  "02112012,23,0.772390    ",
  "03112012,23,0.764040    ",
  "04112012,23,0.755259    ",
  "05112012,23,0.734060    ",
  "06112012,23,0.748574    ",
  "07112012,23,0.766949    ",
  "08112012,23,0.769842    ",
  "09112012,23,0.508916    ",
  "10112012,23,0.084678    ",
  "11112012,23,-0.026953   ",
  "12112012,23,0.028902    ",
  "13112012,23,0.156088    ",
  "14112012,23,0.122295    ",
  "15112012,23,0.019392    ",
  "16112012,23,-0.169461   ",
  "17112012,23,-0.176101   ",
  "18112012,23,-0.177012   ",
  "19112012,23,-0.036819   ",
  "20112012,23,-0.183522   ",
  "21112012,23,-0.130590   ",
  "22112012,23,-0.080360   ",
  "23112012,23,-0.122050   ",
  "24112012,23,-0.145413   ",
  "25112012,23,-0.155407   ",
  "26112012,23,-0.157346   ",
  "27112012,23,-0.173808   ",
  "28112012,23,-0.183500   ",
  "29112012,23,-0.180101   ",
  "30112012,23,-0.176016   ",
  "01122012,23,-0.180731   ",
  "02122012,23,-0.189391   ",
  "03122012,23,-0.179844   ",
  "04122012,23,-0.175133   ",
  "05122012,23,-0.173864   ",
  "06122012,23,-0.164631   ",
  "07122012,23,-0.149067   ",
  "08122012,23,-0.144294   ",
  "09122012,23,-0.137630   ",
  "10122012,23,-0.137132   ",
  "11122012,23,-0.142295   ",
  "12122012,23,-0.141400   ",
  "13122012,23,-0.135970   ",
  "14122012,23,-0.130041   ",
  "15122012,23,-0.128438   ",
  "16122012,23,-0.132093   ",
  "17122012,23,-0.136432   ",
  "18122012,23,-0.133213   ",
  "19122012,23,-0.124260   ",
  "20122012,23,-0.130280   ",
  "21122012,23,-0.129136   ",
  "22122012,23,-0.135866   ",
  "23122012,23,-0.141271   ",
  "24122012,23,-0.138335   ",
  "25122012,23,-0.131582   ",
  "26122012,23,-0.135805   ",
  "27122012,23,-0.129923   ",
  "28122012,23,-0.128358   ",
  "29122012,23,-0.121149   ",
  "30122012,23,-0.117116   ",
  "31122012,23,-0.105243   " ;

 me2012f =
  "17052012  0  0  0  0  5.82829  0  1.23291  0  0  0  0  0  0  0  0  0  0  0  0  0.02  0.76  0  0  1  0  0                        ",
  "16062012  0  0  0  0  0  0  6.72495  0  0  0  0  0  0  0  0  0  0  0  0  0.02  0.76  0  0  1  0  0                              ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                " ;

 me2013t =
  "02042013,3,0.100000     ",
  "01012013,23,-0.105188   ",
  "02012013,23,-0.103553   ",
  "03012013,23,-0.096203   ",
  "04012013,23,-0.095818   ",
  "05012013,23,-0.102792   ",
  "06012013,23,-0.115464   ",
  "07012013,23,-0.117498   ",
  "08012013,23,-0.121575   ",
  "09012013,23,-0.132324   ",
  "10012013,23,-0.123514   ",
  "11012013,23,-0.114553   ",
  "12012013,23,-0.104855   ",
  "13012013,23,-0.096137   ",
  "14012013,23,-0.080427   ",
  "15012013,23,-0.077011   ",
  "16012013,23,-0.088339   ",
  "17012013,23,-0.094770   ",
  "18012013,23,-0.094521   ",
  "19012013,23,-0.091570   ",
  "20012013,23,-0.092431   ",
  "21012013,23,-0.092120   ",
  "22012013,23,-0.094455   ",
  "23012013,23,-0.093355   ",
  "24012013,23,-0.092862   ",
  "25012013,23,-0.102256   ",
  "26012013,23,-0.110296   ",
  "27012013,23,-0.097145   ",
  "28012013,23,-0.093789   ",
  "29012013,23,-0.096220   ",
  "30012013,23,-0.098000   ",
  "31012013,23,-0.104025   ",
  "01022013,23,-0.100365   ",
  "02022013,23,-0.091859   ",
  "03022013,23,-0.091820   ",
  "04022013,23,-0.068068   ",
  "05022013,23,-0.049040   ",
  "06022013,23,-0.032646   ",
  "07022013,23,-0.031332   ",
  "08022013,23,-0.025538   ",
  "09022013,23,-0.005986   ",
  "10022013,23,-0.001515   ",
  "11022013,23,0.013894    ",
  "12022013,23,0.025721    ",
  "13022013,23,0.024643    ",
  "14022013,23,0.034474    ",
  "15022013,23,0.054730    ",
  "16022013,23,0.055661    ",
  "17022013,23,0.068295    ",
  "18022013,23,0.106305    ",
  "19022013,23,0.094682    ",
  "20022013,23,0.088049    ",
  "21022013,23,0.145299    ",
  "22022013,23,0.186817    ",
  "23022013,23,0.210908    ",
  "24022013,23,0.255848    ",
  "25022013,23,0.281931    ",
  "26022013,23,0.298512    ",
  "27022013,23,0.330358    ",
  "28022013,23,0.348840    ",
  "01032013,23,0.347324    ",
  "02032013,23,0.328548    ",
  "03032013,23,0.312812    ",
  "04032013,23,0.336273    ",
  "05032013,23,0.340634    ",
  "06032013,23,0.376265    ",
  "07032013,23,0.376448    ",
  "08032013,23,0.393255    ",
  "09032013,23,0.463192    ",
  "10032013,23,0.479501    ",
  "11032013,23,0.471654    ",
  "12032013,23,0.471901    ",
  "13032013,23,0.485570    ",
  "14032013,23,0.446545    ",
  "15032013,23,0.444010    ",
  "16032013,23,0.458319    ",
  "17032013,23,0.464869    ",
  "18032013,23,0.465602    ",
  "19032013,23,0.460996    ",
  "20032013,23,0.505562    ",
  "21032013,23,0.451140    ",
  "22032013,23,0.478797    ",
  "23032013,23,0.464924    ",
  "24032013,23,0.474848    ",
  "25032013,23,0.473221    ",
  "26032013,23,0.480996    ",
  "27032013,23,0.515415    ",
  "28032013,23,0.552540    ",
  "29032013,23,0.589512    ",
  "30032013,23,0.619625    ",
  "31032013,23,0.647343    ",
  "01042013,23,0.647585    ",
  "02042013,23,0.647151    ",
  "03042013,23,0.653584    ",
  "04042013,23,0.658623    ",
  "05042013,23,0.645382    ",
  "06042013,23,0.633874    ",
  "07042013,23,0.644801    ",
  "08042013,23,0.669568    ",
  "09042013,23,0.657920    ",
  "10042013,23,0.678911    ",
  "11042013,23,0.659926    ",
  "12042013,23,0.625561    ",
  "13042013,23,0.644513    ",
  "14042013,23,0.663896    ",
  "15042013,23,0.681196    ",
  "16042013,23,0.710352    ",
  "17042013,23,0.731206    ",
  "18042013,23,0.739819    ",
  "19042013,23,0.739341    ",
  "20042013,23,0.736240    ",
  "21042013,23,0.741290    ",
  "22042013,23,0.743526    ",
  "23042013,23,0.751122    ",
  "24042013,23,0.757340    ",
  "25042013,23,0.778343    ",
  "26042013,23,0.791821    ",
  "27042013,23,0.791900    ",
  "28042013,23,0.785672    ",
  "29042013,23,0.784476    ",
  "30042013,23,0.794087    ",
  "01052013,23,0.815005    ",
  "02052013,23,0.831629    ",
  "03052013,23,0.829234    ",
  "04052013,23,0.828055    ",
  "05052013,23,0.843075    ",
  "06052013,23,0.860592    ",
  "07052013,23,0.872845    ",
  "08052013,23,0.882160    ",
  "09052013,23,0.894173    ",
  "10052013,23,0.901658    ",
  "11052013,23,0.908570    ",
  "12052013,23,0.915961    ",
  "13052013,23,0.922316    ",
  "14052013,23,0.929967    ",
  "15052013,23,0.932151    ",
  "16052013,23,0.868568    ",
  "17052013,23,0.714139    ",
  "18052013,23,0.014975    ",
  "19052013,23,-0.079328   ",
  "20052013,23,-0.094235   ",
  "21052013,23,-0.103017   ",
  "22052013,23,-0.081129   ",
  "23052013,23,-0.063814   ",
  "24052013,23,-0.056641   ",
  "25052013,23,-0.054548   ",
  "26052013,23,-0.058880   ",
  "27052013,23,-0.064298   ",
  "28052013,23,-0.069846   ",
  "29052013,23,-0.070267   ",
  "30052013,23,-0.071329   ",
  "31052013,23,-0.075015   ",
  "01062013,23,-0.081189   ",
  "02062013,23,-0.084300   ",
  "03062013,23,-0.082190   ",
  "04062013,23,-0.079834   ",
  "05062013,23,-0.076667   ",
  "06062013,23,-0.078008   ",
  "07062013,23,-0.079954   ",
  "08062013,23,-0.080016   ",
  "09062013,23,-0.073465   ",
  "10062013,23,-0.072291   ",
  "11062013,23,-0.076467   ",
  "12062013,23,-0.073368   ",
  "13062013,23,-0.064684   ",
  "14062013,23,-0.064887   ",
  "15062013,23,-0.058088   ",
  "16062013,23,-0.050435   ",
  "17062013,23,-0.047653   ",
  "18062013,23,-0.050093   ",
  "19062013,23,-0.052251   ",
  "20062013,23,-0.057092   ",
  "21062013,23,-0.059490   ",
  "22062013,23,-0.063091   ",
  "23062013,23,-0.064279   ",
  "24062013,23,-0.067234   ",
  "25062013,23,-0.072830   ",
  "26062013,23,-0.073149   ",
  "27062013,23,-0.068875   ",
  "28062013,23,-0.066296   ",
  "29062013,23,-0.064942   ",
  "30062013,23,-0.065940   ",
  "01072013,23,-0.067697   ",
  "02072013,23,-0.075379   ",
  "03072013,23,-0.083744   ",
  "04072013,23,-0.096723   ",
  "05072013,23,-0.086599   ",
  "06072013,23,-0.080598   ",
  "07072013,23,-0.076488   ",
  "08072013,23,-0.071543   ",
  "09072013,23,-0.073884   ",
  "10072013,23,-0.076085   ",
  "11072013,23,-0.072916   ",
  "12072013,23,-0.070307   ",
  "13072013,23,-0.066389   ",
  "14072013,23,-0.066043   ",
  "15072013,23,-0.067405   ",
  "16072013,23,-0.059302   ",
  "17072013,23,-0.057855   ",
  "18072013,23,-0.061112   ",
  "19072013,23,-0.065613   ",
  "20072013,23,-0.071718   ",
  "21072013,23,-0.073204   ",
  "22072013,23,-0.074921   ",
  "23072013,23,-0.087098   ",
  "24072013,23,-0.102617   ",
  "25072013,23,-0.112747   ",
  "26072013,23,-0.085811   ",
  "27072013,23,-0.076384   ",
  "28072013,23,-0.088421   ",
  "29072013,23,-0.098720   ",
  "30072013,23,-0.109016   ",
  "31072013,23,-0.117714   ",
  "01082013,23,-0.124408   ",
  "02082013,23,-0.127241   ",
  "03082013,23,-0.128893   ",
  "04082013,23,-0.131153   ",
  "05082013,23,-0.131759   ",
  "06082013,23,-0.118816   ",
  "07082013,23,-0.105829   ",
  "08082013,23,-0.096503   ",
  "09082013,23,-0.087781   ",
  "10082013,23,-0.078897   ",
  "11082013,23,-0.069504   ",
  "12082013,23,-0.059341   ",
  "13082013,23,-0.049862   ",
  "14082013,23,-0.036828   ",
  "15082013,23,-0.024941   ",
  "16082013,23,-0.015278   ",
  "17082013,23,-0.006088   ",
  "18082013,23,0.001836    ",
  "19082013,23,0.011593    ",
  "20082013,23,0.026907    ",
  "21082013,23,0.050478    ",
  "22082013,23,0.068168    ",
  "23082013,23,0.090623    ",
  "24082013,23,0.163227    ",
  "25082013,23,0.230120    ",
  "26082013,23,0.285550    ",
  "27082013,23,0.327791    ",
  "28082013,23,0.391538    ",
  "29082013,23,0.446922    ",
  "30082013,23,0.480486    ",
  "31082013,23,0.522086    ",
  "01092013,23,0.569956    ",
  "02092013,23,0.619773    ",
  "03092013,23,0.664790    ",
  "04092013,23,0.710429    ",
  "05092013,23,0.750062    ",
  "06092013,23,0.786872    ",
  "07092013,23,0.818696    ",
  "08092013,23,0.849959    ",
  "09092013,23,0.876686    ",
  "10092013,23,0.912391    ",
  "11092013,23,0.945019    ",
  "12092013,23,0.962726    ",
  "13092013,23,0.974196    ",
  "14092013,23,0.936817    ",
  "15092013,23,0.928156    ",
  "16092013,23,0.928290    ",
  "17092013,23,0.928173    ",
  "18092013,23,0.921133    ",
  "19092013,23,0.908039    ",
  "20092013,23,0.931051    ",
  "21092013,23,0.926183    ",
  "22092013,23,0.929876    ",
  "23092013,23,0.930423    ",
  "24092013,23,0.888023    ",
  "25092013,23,0.825231    ",
  "26092013,23,0.919598    ",
  "27092013,23,0.870371    ",
  "28092013,23,0.529682    ",
  "29092013,23,0.848615    ",
  "30092013,23,0.847379    ",
  "01102013,23,0.710992    ",
  "02102013,23,0.449723    ",
  "03102013,23,0.281361    ",
  "04102013,23,-0.032914   ",
  "05102013,23,-0.014431   ",
  "06102013,23,-0.032979   ",
  "07102013,23,-0.120903   ",
  "08102013,23,-0.112935   ",
  "09102013,23,-0.154888   ",
  "10102013,23,-0.186871   ",
  "11102013,23,-0.189205   ",
  "12102013,23,-0.204519   ",
  "13102013,23,-0.210655   ",
  "14102013,23,-0.206905   ",
  "15102013,23,-0.207190   ",
  "16102013,23,-0.205377   ",
  "17102013,23,-0.166590   ",
  "18102013,23,-0.203765   ",
  "19102013,23,-0.218223   ",
  "20102013,23,-0.226300   ",
  "21102013,23,-0.233622   ",
  "22102013,23,-0.240325   ",
  "23102013,23,-0.247360   ",
  "24102013,23,-0.253756   ",
  "25102013,23,-0.256827   ",
  "26102013,23,-0.262547   ",
  "27102013,23,-0.263413   ",
  "28102013,23,-0.227060   ",
  "29102013,23,-0.224621   ",
  "30102013,23,-0.223736   ",
  "31102013,23,-0.220973   ",
  "01112013,23,-0.215143   ",
  "02112013,23,-0.212969   ",
  "03112013,23,-0.208469   ",
  "04112013,23,-0.207997   ",
  "05112013,23,-0.211845   ",
  "06112013,23,-0.207559   ",
  "07112013,23,-0.192620   ",
  "08112013,23,-0.173664   ",
  "09112013,23,-0.161369   ",
  "10112013,23,-0.170597   ",
  "11112013,23,-0.172260   ",
  "12112013,23,-0.169320   ",
  "13112013,23,-0.169092   ",
  "14112013,23,-0.166245   ",
  "15112013,23,-0.141001   ",
  "16112013,23,-0.143703   ",
  "17112013,23,-0.142593   ",
  "18112013,23,-0.146249   ",
  "19112013,23,-0.148179   ",
  "20112013,23,-0.147424   ",
  "21112013,23,-0.144511   ",
  "22112013,23,-0.142032   ",
  "23112013,23,-0.137669   ",
  "24112013,23,-0.134108   ",
  "25112013,23,-0.131563   ",
  "26112013,23,-0.128621   ",
  "27112013,23,-0.126016   ",
  "28112013,23,-0.120739   ",
  "29112013,23,-0.110122   ",
  "30112013,23,-0.096163   ",
  "01122013,23,-0.086271   ",
  "02122013,23,-0.081861   ",
  "03122013,23,-0.105702   ",
  "04122013,23,-0.086030   ",
  "05122013,23,-0.075327   ",
  "06122013,23,-0.071655   ",
  "07122013,23,-0.096785   ",
  "08122013,23,-0.088485   ",
  "09122013,23,-0.081868   ",
  "10122013,23,-0.077718   ",
  "11122013,23,-0.074619   ",
  "12122013,23,-0.071334   ",
  "13122013,23,-0.070747   ",
  "14122013,23,-0.069470   ",
  "15122013,23,-0.068777   ",
  "16122013,23,-0.067980   ",
  "17122013,23,-0.067186   ",
  "18122013,23,-0.067137   ",
  "19122013,23,-0.093468   ",
  "20122013,23,-0.099831   ",
  "21122013,23,-0.097427   ",
  "22122013,23,-0.095328   ",
  "23122013,23,-0.094270   ",
  "24122013,23,-0.094231   ",
  "25122013,23,-0.093877   ",
  "26122013,23,-0.093830   ",
  "27122013,23,-0.094077   ",
  "28122013,23,-0.095095   ",
  "29122013,23,-0.092601   ",
  "30122013,23,-0.093590   ",
  "31122013,23,-0.095415   ",
  "                        " ;

 me2013f =
  "02052013  0  0  0  0  1.68124  0  1.68124  0  0  0  0  0  0  0  0  0  0  0  0  0.02  0.76  0  0  1  0  0                        ",
  "16062013  0  0  0  0  0  0  6.72495  0  0  0  0  0  0  0  0  0  0  0  0  0.02  0.76  0  0  1  0  0                              ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                " ;

 me2014t =
  "28042014,3,0.100000     ",
  "01012014,23,-0.097365   ",
  "02012014,23,-0.099113   ",
  "03012014,23,-0.101202   ",
  "04012014,23,-0.101103   ",
  "05012014,23,-0.099082   ",
  "06012014,23,-0.099462   ",
  "07012014,23,-0.101188   ",
  "08012014,23,-0.103211   ",
  "09012014,23,-0.106179   ",
  "10012014,23,-0.102286   ",
  "11012014,23,-0.105439   ",
  "12012014,23,-0.103891   ",
  "13012014,23,-0.098090   ",
  "14012014,23,-0.098537   ",
  "15012014,23,-0.099233   ",
  "16012014,23,-0.099584   ",
  "17012014,23,-0.099532   ",
  "18012014,23,-0.100201   ",
  "19012014,23,-0.099935   ",
  "20012014,23,-0.098953   ",
  "21012014,23,-0.098400   ",
  "22012014,23,-0.099579   ",
  "23012014,23,-0.100641   ",
  "24012014,23,-0.099864   ",
  "25012014,23,-0.098464   ",
  "26012014,23,-0.094913   ",
  "27012014,23,-0.087505   ",
  "28012014,23,-0.080479   ",
  "29012014,23,-0.075292   ",
  "30012014,23,-0.073201   ",
  "31012014,23,-0.071781   ",
  "01022014,23,-0.074535   ",
  "02022014,23,-0.065642   ",
  "03022014,23,-0.057452   ",
  "04022014,23,-0.043045   ",
  "05022014,23,-0.033195   ",
  "06022014,23,-0.032228   ",
  "07022014,23,-0.030036   ",
  "08022014,23,-0.084121   ",
  "09022014,23,-0.121393   ",
  "10022014,23,-0.135368   ",
  "11022014,23,-0.144916   ",
  "12022014,23,-0.180727   ",
  "13022014,23,-0.170510   ",
  "14022014,23,-0.143844   ",
  "15022014,23,-0.111070   ",
  "16022014,23,-0.083696   ",
  "17022014,23,-0.061274   ",
  "18022014,23,-0.043017   ",
  "19022014,23,-0.028812   ",
  "20022014,23,-0.016734   ",
  "21022014,23,-0.008564   ",
  "22022014,23,0.003147    ",
  "23022014,23,0.012214    ",
  "24022014,23,0.018989    ",
  "25022014,23,0.027895    ",
  "26022014,23,0.020099    ",
  "27022014,23,0.003789    ",
  "28022014,23,-0.008054   ",
  "01032014,23,0.001269    ",
  "02032014,23,0.012707    ",
  "03032014,23,0.015098    ",
  "04032014,23,0.013245    ",
  "05032014,23,0.013391    ",
  "06032014,23,0.016954    ",
  "07032014,23,0.030694    ",
  "08032014,23,0.051565    ",
  "09032014,23,0.056286    ",
  "10032014,23,0.082128    ",
  "11032014,23,0.136320    ",
  "12032014,23,0.202226    ",
  "13032014,23,0.244569    ",
  "14032014,23,0.288615    ",
  "15032014,23,0.316256    ",
  "16032014,23,0.329635    ",
  "17032014,23,0.342400    ",
  "18032014,23,0.376479    ",
  "19032014,23,0.419725    ",
  "20032014,23,0.430090    ",
  "21032014,23,0.445888    ",
  "22032014,23,0.480230    ",
  "23032014,23,0.500995    ",
  "24032014,23,0.508752    ",
  "25032014,23,0.507524    ",
  "26032014,23,0.492314    ",
  "27032014,23,0.486744    ",
  "28032014,23,0.488565    ",
  "29032014,23,0.449219    ",
  "30032014,23,0.402268    ",
  "31032014,23,0.376194    ",
  "01042014,23,0.273110    ",
  "02042014,23,0.193651    ",
  "03042014,23,0.225491    ",
  "04042014,23,0.218566    ",
  "05042014,23,0.229880    ",
  "06042014,23,0.263686    ",
  "07042014,23,0.286475    ",
  "08042014,23,0.303623    ",
  "09042014,23,0.322575    ",
  "10042014,23,0.341415    ",
  "11042014,23,0.356149    ",
  "12042014,23,0.383502    ",
  "13042014,23,0.424471    ",
  "14042014,23,0.453199    ",
  "15042014,23,0.459486    ",
  "16042014,23,0.476089    ",
  "17042014,23,0.422953    ",
  "18042014,23,0.427304    ",
  "19042014,23,0.427298    ",
  "20042014,23,0.453062    ",
  "21042014,23,0.436267    ",
  "22042014,23,0.447195    ",
  "23042014,23,0.436017    ",
  "24042014,23,0.443658    ",
  "25042014,23,0.446092    ",
  "26042014,23,0.437886    ",
  "27042014,23,0.453551    ",
  "28042014,23,0.455547    ",
  "29042014,23,0.457648    ",
  "30042014,23,0.473587    ",
  "01052014,23,0.464667    ",
  "02052014,23,0.432193    ",
  "03052014,23,0.436919    ",
  "04052014,23,0.453502    ",
  "05052014,23,0.460116    ",
  "06052014,23,0.461116    ",
  "07052014,23,0.481282    ",
  "08052014,23,0.501158    ",
  "09052014,23,0.511365    ",
  "10052014,23,0.511514    ",
  "11052014,23,0.517603    ",
  "12052014,23,0.526430    ",
  "13052014,23,0.533765    ",
  "14052014,23,0.533208    ",
  "15052014,23,0.533922    ",
  "16052014,23,0.535073    ",
  "17052014,23,0.540949    ",
  "18052014,23,0.552760    ",
  "19052014,23,0.562367    ",
  "20052014,23,0.576231    ",
  "21052014,23,0.580631    ",
  "22052014,23,0.589159    ",
  "23052014,23,0.596209    ",
  "24052014,23,0.604458    ",
  "25052014,23,0.615325    ",
  "26052014,23,0.630779    ",
  "27052014,23,0.648549    ",
  "28052014,23,0.651630    ",
  "29052014,23,0.648493    ",
  "30052014,23,0.648478    ",
  "31052014,23,0.648583    ",
  "01062014,23,0.648611    ",
  "02062014,23,0.648341    ",
  "03062014,23,0.648537    ",
  "04062014,23,0.648554    ",
  "05062014,23,0.648488    ",
  "06062014,23,0.648432    ",
  "07062014,23,0.648479    ",
  "08062014,23,0.647387    ",
  "09062014,23,0.400651    ",
  "10062014,23,-0.170893   ",
  "11062014,23,-0.226066   ",
  "12062014,23,-0.238555   ",
  "13062014,23,-0.240957   ",
  "14062014,23,-0.238816   ",
  "15062014,23,-0.239385   ",
  "16062014,23,-0.235315   ",
  "17062014,23,-0.207528   ",
  "18062014,23,-0.211565   ",
  "19062014,23,-0.215953   ",
  "20062014,23,-0.218124   ",
  "21062014,23,-0.219983   ",
  "22062014,23,-0.222187   ",
  "23062014,23,-0.224690   ",
  "24062014,23,-0.223352   ",
  "25062014,23,-0.223680   ",
  "26062014,23,-0.222350   ",
  "27062014,23,-0.222862   ",
  "28062014,23,-0.228789   ",
  "29062014,23,-0.233799   ",
  "30062014,23,-0.239514   ",
  "01072014,23,-0.243805   ",
  "02072014,23,-0.244883   ",
  "03072014,23,-0.246739   ",
  "04072014,23,-0.248382   ",
  "05072014,23,-0.250011   ",
  "06072014,23,-0.253534   ",
  "07072014,23,-0.259604   ",
  "08072014,23,-0.249644   ",
  "09072014,23,-0.230338   ",
  "10072014,23,-0.230062   ",
  "11072014,23,-0.228902   ",
  "12072014,23,-0.227951   ",
  "13072014,23,-0.224340   ",
  "14072014,23,-0.221444   ",
  "15072014,23,-0.216566   ",
  "16072014,23,-0.213750   ",
  "17072014,23,-0.217031   ",
  "18072014,23,-0.218066   ",
  "19072014,23,-0.216055   ",
  "20072014,23,-0.214183   ",
  "21072014,23,-0.207060   ",
  "22072014,23,-0.201845   ",
  "23072014,23,-0.192838   ",
  "24072014,23,-0.184524   ",
  "25072014,23,-0.189392   ",
  "26072014,23,-0.191041   ",
  "27072014,23,-0.190216   ",
  "28072014,23,-0.189439   ",
  "29072014,23,-0.190054   ",
  "30072014,23,-0.193473   ",
  "31072014,23,-0.204855   ",
  "01082014,23,-0.208346   ",
  "02082014,23,-0.205332   ",
  "03082014,23,-0.202497   ",
  "04082014,23,-0.199898   ",
  "05082014,23,-0.195687   ",
  "06082014,23,-0.193134   ",
  "07082014,23,-0.192783   ",
  "08082014,23,-0.194768   ",
  "09082014,23,-0.195395   ",
  "10082014,23,-0.191450   ",
  "11082014,23,-0.180800   ",
  "12082014,23,-0.177889   ",
  "13082014,23,-0.169342   ",
  "14082014,23,-0.158682   ",
  "15082014,23,-0.149746   ",
  "16082014,23,-0.141985   ",
  "17082014,23,-0.134939   ",
  "18082014,23,-0.131295   ",
  "19082014,23,-0.153737   ",
  "20082014,23,-0.176009   ",
  "21082014,23,-0.158627   ",
  "22082014,23,-0.148026   ",
  "23082014,23,-0.134543   ",
  "24082014,23,-0.119095   ",
  "25082014,23,-0.067138   ",
  "26082014,23,-0.007570   ",
  "27082014,23,0.055528    ",
  "28082014,23,0.108440    ",
  "29082014,23,0.159232    ",
  "30082014,23,0.216424    ",
  "31082014,23,0.274418    ",
  "01092014,23,0.313358    ",
  "02092014,23,0.350857    ",
  "03092014,23,0.394002    ",
  "04092014,23,0.437469    ",
  "05092014,23,0.493837    ",
  "06092014,23,0.532894    ",
  "07092014,23,0.563049    ",
  "08092014,23,0.600169    ",
  "09092014,23,0.635610    ",
  "10092014,23,0.654643    ",
  "11092014,23,0.650837    ",
  "12092014,23,0.648169    ",
  "13092014,23,0.648172    ",
  "14092014,23,0.648179    ",
  "15092014,23,0.648195    ",
  "16092014,23,0.648209    ",
  "17092014,23,0.648213    ",
  "18092014,23,0.648228    ",
  "19092014,23,0.648240    ",
  "20092014,23,0.648256    ",
  "21092014,23,0.648291    ",
  "22092014,23,0.648280    ",
  "23092014,23,0.648282    ",
  "24092014,23,0.648294    ",
  "25092014,23,0.648300    ",
  "26092014,23,0.648317    ",
  "27092014,23,0.648315    ",
  "28092014,23,0.648330    ",
  "29092014,23,0.648331    ",
  "30092014,23,0.648308    ",
  "01102014,23,0.648257    ",
  "02102014,23,0.648310    ",
  "03102014,23,0.648311    ",
  "04102014,23,0.648311    ",
  "05102014,23,0.648295    ",
  "06102014,23,0.648295    ",
  "07102014,23,0.648273    ",
  "08102014,23,0.648702    ",
  "09102014,23,0.648287    ",
  "10102014,23,0.648311    ",
  "11102014,23,0.647415    ",
  "12102014,23,0.569023    ",
  "13102014,23,0.456442    ",
  "14102014,23,0.515997    ",
  "15102014,23,0.427173    ",
  "16102014,23,0.484534    ",
  "17102014,23,0.426428    ",
  "18102014,23,0.229089    ",
  "19102014,23,0.097926    ",
  "20102014,23,-0.011416   ",
  "21102014,23,-0.018505   ",
  "22102014,23,-0.009049   ",
  "23102014,23,0.062614    ",
  "24102014,23,0.204880    ",
  "25102014,23,-0.045860   ",
  "26102014,23,0.019198    ",
  "27102014,23,0.052994    ",
  "28102014,23,-0.013571   ",
  "29102014,23,0.006512    ",
  "30102014,23,0.279468    ",
  "31102014,23,-0.087503   ",
  "01112014,23,-0.082375   ",
  "02112014,23,-0.076638   ",
  "03112014,23,-0.070798   ",
  "04112014,23,-0.067799   ",
  "05112014,23,-0.066717   ",
  "06112014,23,-0.062354   ",
  "07112014,23,-0.061853   ",
  "08112014,23,-0.060361   ",
  "09112014,23,-0.062183   ",
  "10112014,23,-0.061577   ",
  "11112014,23,-0.065932   ",
  "12112014,23,-0.074061   ",
  "13112014,23,-0.085299   ",
  "14112014,23,-0.096439   ",
  "15112014,23,-0.100297   ",
  "16112014,23,-0.104601   ",
  "17112014,23,-0.110235   ",
  "18112014,23,-0.113591   ",
  "19112014,23,-0.118425   ",
  "20112014,23,-0.127076   ",
  "21112014,23,-0.134604   ",
  "22112014,23,-0.148168   ",
  "23112014,23,-0.161679   ",
  "24112014,23,-0.162845   ",
  "25112014,23,-0.161054   ",
  "26112014,23,-0.162631   ",
  "27112014,23,-0.164601   ",
  "28112014,23,-0.164395   ",
  "29112014,23,-0.159000   ",
  "30112014,23,-0.152099   ",
  "01122014,23,-0.153802   ",
  "02122014,23,-0.174882   ",
  "03122014,23,-0.206354   ",
  "04122014,23,-0.230096   ",
  "05122014,23,-0.232336   ",
  "06122014,23,-0.226910   ",
  "07122014,23,-0.217348   ",
  "08122014,23,-0.200908   ",
  "09122014,23,-0.183551   ",
  "10122014,23,-0.197568   ",
  "11122014,23,-0.220968   ",
  "12122014,23,-0.203862   ",
  "13122014,23,-0.217750   ",
  "14122014,23,-0.222650   ",
  "15122014,23,-0.227575   ",
  "16122014,23,-0.235946   ",
  "17122014,23,-0.248069   ",
  "18122014,23,-0.248221   ",
  "19122014,23,-0.243210   ",
  "20122014,23,-0.244160   ",
  "21122014,23,-0.242204   ",
  "22122014,23,-0.232359   ",
  "23122014,23,-0.212361   ",
  "24122014,23,-0.199363   ",
  "25122014,23,-0.171580   ",
  "26122014,23,-0.138905   ",
  "27122014,23,-0.114451   ",
  "28122014,23,-0.105276   ",
  "29122014,23,-0.099440   ",
  "30122014,23,-0.092068   ",
  "31122014,23,-0.082664   ",
  "                        " ;

 me2014f =
  "05062014  0  0  0  0  2.52186  0  2.52186  0  0  0  0  0  0  0  0  0  0  0  0  0.02  0.76  0  0  1  0  0                        ",
  "16062014  0  0  0  0  0  0  6.72495  0  0  0  0  0  0  0  0  0  0  0  0  0.02  0.76  0  0  1  0  0                              ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                " ;

 me2015t =
  "16042015,3,0.100000     ",
  "01012015,23,-0.065728   ",
  "02012015,23,-0.059226   ",
  "03012015,23,-0.049022   ",
  "04012015,23,-0.042687   ",
  "05012015,23,-0.041823   ",
  "06012015,23,-0.038964   ",
  "07012015,23,-0.037946   ",
  "08012015,23,-0.036579   ",
  "09012015,23,-0.034676   ",
  "10012015,23,-0.033566   ",
  "11012015,23,-0.030336   ",
  "12012015,23,-0.031069   ",
  "13012015,23,-0.032692   ",
  "14012015,23,-0.029984   ",
  "15012015,23,-0.032241   ",
  "16012015,23,-0.033077   ",
  "17012015,23,-0.032614   ",
  "18012015,23,-0.029685   ",
  "19012015,23,-0.030606   ",
  "20012015,23,-0.027457   ",
  "21012015,23,-0.019764   ",
  "22012015,23,-0.014186   ",
  "23012015,23,-0.015248   ",
  "24012015,23,-0.015065   ",
  "25012015,23,-0.015233   ",
  "26012015,23,-0.015481   ",
  "27012015,23,-0.006885   ",
  "28012015,23,-0.011720   ",
  "29012015,23,-0.010718   ",
  "30012015,23,-0.009592   ",
  "31012015,23,0.003218    ",
  "01022015,23,0.017159    ",
  "02022015,23,0.036638    ",
  "03022015,23,0.054091    ",
  "04022015,23,0.063560    ",
  "05022015,23,0.070205    ",
  "06022015,23,0.070922    ",
  "07022015,23,0.070829    ",
  "08022015,23,0.060917    ",
  "09022015,23,0.076581    ",
  "10022015,23,0.079288    ",
  "11022015,23,0.087929    ",
  "12022015,23,0.091185    ",
  "13022015,23,0.093491    ",
  "14022015,23,0.098909    ",
  "15022015,23,0.105843    ",
  "16022015,23,0.114950    ",
  "17022015,23,0.136766    ",
  "18022015,23,0.152260    ",
  "19022015,23,0.149811    ",
  "20022015,23,0.146430    ",
  "21022015,23,0.162250    ",
  "22022015,23,0.197832    ",
  "23022015,23,0.291266    ",
  "24022015,23,0.345934    ",
  "25022015,23,0.340017    ",
  "26022015,23,0.333197    ",
  "27022015,23,0.355823    ",
  "28022015,23,0.402296    ",
  "01032015,23,0.428324    ",
  "02032015,23,0.425302    ",
  "03032015,23,0.453434    ",
  "04032015,23,0.483884    ",
  "08052015,23,0.021766    ",
  "09052015,23,0.051896    ",
  "10052015,23,0.067361    ",
  "11052015,23,0.100407    ",
  "12052015,23,0.179104    ",
  "13052015,23,0.246563    ",
  "14052015,23,0.273399    ",
  "15052015,23,0.317144    ",
  "16052015,23,0.373288    ",
  "17052015,23,0.414938    ",
  "18052015,23,0.452263    ",
  "19052015,23,0.477888    ",
  "20052015,23,0.493878    ",
  "21052015,23,0.524912    ",
  "22052015,23,0.561852    ",
  "23052015,23,0.590136    ",
  "24052015,23,0.604135    ",
  "25052015,23,0.634607    ",
  "26052015,23,0.669600    ",
  "27052015,23,0.696124    ",
  "28052015,23,0.717851    ",
  "29052015,23,0.738105    ",
  "30052015,23,0.756984    ",
  "31052015,23,0.742728    ",
  "01062015,23,0.681421    ",
  "02062015,23,0.585586    ",
  "03062015,23,0.431183    ",
  "04062015,23,0.293739    ",
  "05062015,23,0.221564    ",
  "06062015,23,0.156694    ",
  "07062015,23,0.027536    ",
  "08062015,23,-0.011515   ",
  "09062015,23,-0.035994   ",
  "10062015,23,-0.039037   ",
  "11062015,23,-0.056971   ",
  "12062015,23,-0.056263   ",
  "13062015,23,-0.042628   ",
  "14062015,23,-0.030746   ",
  "15062015,23,-0.019166   ",
  "16062015,23,-0.008821   ",
  "17062015,23,-0.000508   ",
  "18062015,23,0.000627    ",
  "19062015,23,0.008162    ",
  "20062015,23,0.027269    ",
  "21062015,23,0.047411    ",
  "22062015,23,0.082193    ",
  "23062015,23,0.104153    ",
  "24062015,23,0.026722    ",
  "25062015,23,-0.009224   ",
  "26062015,23,-0.028573   ",
  "27062015,23,-0.048255   ",
  "28062015,23,-0.070321   ",
  "29062015,23,-0.092272   ",
  "30062015,23,-0.112811   ",
  "01072015,23,-0.129699   ",
  "02072015,23,-0.143284   ",
  "03072015,23,-0.154871   ",
  "04072015,23,-0.163982   ",
  "05072015,23,-0.169244   ",
  "06072015,23,-0.173219   ",
  "07072015,23,-0.179553   ",
  "08072015,23,-0.185527   ",
  "09072015,23,-0.190836   ",
  "10072015,23,-0.197891   ",
  "11072015,23,-0.204973   ",
  "12072015,23,-0.203340   ",
  "13072015,23,-0.206840   ",
  "14072015,23,-0.211361   ",
  "15072015,23,-0.214565   ",
  "16072015,23,-0.223702   ",
  "17072015,23,-0.240827   ",
  "18072015,23,-0.254164   ",
  "19072015,23,-0.264410   ",
  "20072015,23,-0.284423   ",
  "21072015,23,-0.263999   ",
  "22072015,23,-0.235912   ",
  "23072015,23,-0.229839   ",
  "24072015,23,-0.218864   ",
  "25072015,23,-0.215586   ",
  "26072015,23,-0.223313   ",
  "27072015,23,-0.222908   ",
  "28072015,23,-0.225828   ",
  "29072015,23,-0.237862   ",
  "30072015,23,-0.228958   ",
  "31072015,23,-0.241792   ",
  "01082015,23,-0.242832   ",
  "02082015,23,-0.243625   ",
  "03082015,23,-0.218022   ",
  "04082015,23,-0.196749   ",
  "05082015,23,-0.173862   ",
  "06082015,23,-0.147440   ",
  "07082015,23,-0.123435   ",
  "08082015,23,-0.091480   ",
  "09082015,23,-0.057910   ",
  "10082015,23,-0.027194   ",
  "11082015,23,-0.003984   ",
  "12082015,23,0.012902    ",
  "13082015,23,0.029336    ",
  "14082015,23,0.075828    ",
  "15082015,23,0.134701    ",
  "16082015,23,0.190585    ",
  "17082015,23,0.246491    ",
  "18082015,23,0.319962    ",
  "19082015,23,0.376181    ",
  "20082015,23,0.420894    ",
  "21082015,23,0.470230    ",
  "22082015,23,0.507842    ",
  "23082015,23,0.551131    ",
  "24082015,23,0.595378    ",
  "25082015,23,0.618715    ",
  "26082015,23,0.637704    ",
  "27082015,23,0.637700    ",
  "28082015,23,0.637710    ",
  "29082015,23,0.637704    ",
  "30082015,23,0.637698    ",
  "31082015,23,0.637730    ",
  "01092015,23,0.637739    ",
  "02092015,23,0.637715    ",
  "03092015,23,0.637731    ",
  "04092015,23,0.637745    ",
  "05092015,23,0.637777    ",
  "06092015,23,0.637779    ",
  "07092015,23,0.637775    ",
  "08092015,23,0.637777    ",
  "09092015,23,0.637771    ",
  "10092015,23,0.637778    ",
  "11092015,23,0.637774    ",
  "12092015,23,0.637768    ",
  "13092015,23,0.637772    ",
  "14092015,23,0.637749    ",
  "15092015,23,0.637750    ",
  "16092015,23,0.637759    ",
  "17092015,23,0.647551    ",
  "18092015,23,0.692683    ",
  "19092015,23,0.674649    ",
  "20092015,23,0.658446    ",
  "21092015,23,0.679604    ",
  "22092015,23,0.775014    ",
  "23092015,23,0.786067    ",
  "24092015,23,0.788549    ",
  "25092015,23,0.813747    ",
  "26092015,23,0.818223    ",
  "27092015,23,0.821919    ",
  "28092015,23,0.821497    ",
  "29092015,23,0.816740    ",
  "30092015,23,0.817745    ",
  "01102015,23,0.817697    ",
  "02102015,23,0.817622    ",
  "03102015,23,0.817714    ",
  "04102015,23,0.817740    ",
  "05102015,23,0.817911    ",
  "06102015,23,0.817692    ",
  "07102015,23,0.817793    ",
  "08102015,23,0.816686    ",
  "09102015,23,0.782676    ",
  "10102015,23,0.769573    ",
  "11102015,23,0.728439    ",
  "12102015,23,0.719680    ",
  "13102015,23,0.723916    ",
  "14102015,23,0.755886    ",
  "15102015,23,0.726833    ",
  "16102015,23,0.759620    ",
  "17102015,23,0.686477    ",
  "18102015,23,0.673758    ",
  "19102015,23,0.675448    ",
  "20102015,23,0.710723    ",
  "21102015,23,0.663245    ",
  "22102015,23,0.667339    ",
  "23102015,23,0.655977    ",
  "24102015,23,0.647253    ",
  "25102015,23,0.691652    ",
  "26102015,23,0.658201    ",
  "27102015,23,0.653368    ",
  "28102015,23,0.685968    ",
  "29102015,23,0.678493    ",
  "30102015,23,0.644090    ",
  "31102015,23,0.638923    ",
  "01112015,23,0.434702    ",
  "02112015,23,0.273569    ",
  "03112015,23,0.182388    ",
  "04112015,23,-0.007701   ",
  "05112015,23,-0.166128   ",
  "06112015,23,-0.074649   ",
  "07112015,23,-0.042705   ",
  "08112015,23,-0.008450   ",
  "09112015,23,-0.036611   ",
  "10112015,23,-0.194798   ",
  "11112015,23,-0.309694   ",
  "12112015,23,-0.190304   ",
  "13112015,23,-0.115253   ",
  "14112015,23,-0.062878   ",
  "15112015,23,-0.066381   ",
  "16112015,23,-0.338201   ",
  "17112015,23,-0.349720   ",
  "18112015,23,-0.241546   ",
  "19112015,23,-0.158868   ",
  "20112015,23,-0.105541   ",
  "21112015,23,-0.084564   ",
  "22112015,23,-0.071088   ",
  "23112015,23,-0.043579   ",
  "24112015,23,-0.047354   ",
  "25112015,23,-0.151532   ",
  "26112015,23,-0.294560   ",
  "27112015,23,-0.360716   ",
  "28112015,23,-0.379969   ",
  "29112015,23,-0.381425   ",
  "30112015,23,-0.382504   ",
  "01122015,23,-0.337857   ",
  "02122015,23,-0.209124   ",
  "03122015,23,-0.130226   ",
  "04122015,23,-0.221873   ",
  "05122015,23,-0.236188   ",
  "06122015,23,-0.178888   ",
  "07122015,23,-0.135007   ",
  "08122015,23,-0.109054   ",
  "09122015,23,-0.033843   ",
  "10122015,23,0.050080    ",
  "11122015,23,0.001788    ",
  "12122015,23,-0.178420   ",
  "13122015,23,-0.081251   ",
  "14122015,23,-0.229912   ",
  "15122015,23,-0.163126   ",
  "16122015,23,-0.174275   ",
  "17122015,23,-0.156864   ",
  "18122015,23,-0.057074   ",
  "19122015,23,-0.014548   ",
  "20122015,23,-0.156532   ",
  "21122015,23,0.006158    ",
  "22122015,23,0.057873    ",
  "23122015,23,-0.061766   ",
  "24122015,23,-0.025580   ",
  "25122015,23,-0.211300   ",
  "26122015,23,-0.237165   ",
  "27122015,23,-0.161176   ",
  "28122015,23,0.003022    ",
  "29122015,23,-0.017772   ",
  "30122015,23,-0.114237   ",
  "31122015,23,-0.057911   ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        ",
  "                        " ;

 me2015f =
  "31052015  0  0  0  0  1.68124  0  1.68124  0  0  0  0  0  0  0  0  0  0  0  0  0.02  0.76  0  0  1  0  0                        ",
  "16062015  0  0  0  0  0  0  6.72495  0  0  0  0  0  0  0  0  0  0  0  0  0.02  0.76  0  0  1  0  0                              ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                " ;

 me2016t =
  "16042016,3,0.100000     ",
  "01012016,23,-0.054502   ",
  "02012016,23,-0.003858   ",
  "03012016,23,0.098110    ",
  "04012016,23,0.176105    ",
  "05012016,23,0.202651    ",
  "06012016,23,0.208754    ",
  "07012016,23,0.083793    ",
  "08012016,23,0.014636    ",
  "09012016,23,0.032548    ",
  "10012016,23,0.028895    ",
  "11012016,23,-0.000439   ",
  "12012016,23,0.043108    ",
  "13012016,23,0.052578    ",
  "14012016,23,0.030710    ",
  "15012016,23,0.042570    ",
  "16012016,23,0.076261    ",
  "17012016,23,0.084124    ",
  "18012016,23,0.072650    ",
  "19012016,23,0.058562    ",
  "20012016,23,0.034524    ",
  "21012016,23,0.069663    ",
  "22012016,23,0.109479    ",
  "23012016,23,0.071428    ",
  "24012016,23,-0.049004   ",
  "25012016,23,-0.003478   ",
  "26012016,23,-0.006296   ",
  "27012016,23,0.007573    ",
  "28012016,23,0.034123    ",
  "29012016,23,0.112823    ",
  "30012016,23,0.142166    ",
  "31012016,23,0.190772    ",
  "01022016,23,-0.093029   ",
  "02022016,23,-0.067790   ",
  "03022016,23,-0.095000   ",
  "04022016,23,-0.034182   ",
  "05022016,23,0.000447    ",
  "06022016,23,0.028592    ",
  "07022016,23,0.106669    ",
  "08022016,23,0.146576    ",
  "09022016,23,0.168065    ",
  "10022016,23,0.176581    ",
  "11022016,23,0.208965    ",
  "12022016,23,0.207238    ",
  "13022016,23,0.223640    ",
  "14022016,23,0.270928    ",
  "15022016,23,0.367639    ",
  "16022016,23,0.447899    ",
  "17022016,23,0.558686    ",
  "18022016,23,0.400346    ",
  "19022016,23,0.328083    ",
  "20022016,23,0.301236    ",
  "21022016,23,0.290536    ",
  "22022016,23,0.329930    ",
  "23022016,23,0.383002    ",
  "24022016,23,0.389324    ",
  "25022016,23,0.427174    ",
  "26022016,23,0.462040    ",
  "27022016,23,0.481399    ",
  "28022016,23,0.498310    ",
  "29022016,23,0.533654    ",
  "01032016,23,0.588924    ",
  "02032016,23,0.644076    ",
  "03032016,23,0.672422    ",
  "04032016,23,0.663198    ",
  "05032016,23,0.582212    ",
  "06032016,23,0.463841    ",
  "07032016,23,0.446110    ",
  "08032016,23,0.335487    ",
  "09032016,23,0.395385    ",
  "10032016,23,0.449146    ",
  "11032016,23,0.480451    ",
  "12032016,23,0.338236    ",
  "13032016,23,0.400986    ",
  "14032016,23,0.343721    ",
  "15032016,23,0.344889    ",
  "16032016,23,0.397875    ",
  "17032016,23,0.463298    ",
  "18032016,23,0.475675    ",
  "19032016,23,0.486731    ",
  "20032016,23,0.474769    ",
  "21032016,23,0.465029    ",
  "22032016,23,0.412907    ",
  "23032016,23,0.439947    ",
  "24032016,23,0.533800    ",
  "25032016,23,0.646312    ",
  "26032016,23,0.729209    ",
  "27032016,23,0.763305    ",
  "28032016,23,0.761759    ",
  "29032016,23,0.807269    ",
  "30032016,23,0.846997    ",
  "31032016,23,0.833242    ",
  "01042016,23,0.832154    ",
  "02042016,23,0.845023    ",
  "03042016,23,0.877130    ",
  "04042016,23,0.877159    ",
  "05042016,23,0.878941    ",
  "06042016,23,0.939765    ",
  "07042016,23,0.981690    ",
  "08042016,23,0.988961    ",
  "09042016,23,0.939328    ",
  "10042016,23,0.910005    ",
  "11042016,23,0.903371    ",
  "12042016,23,0.854642    ",
  "13042016,23,0.927734    ",
  "14042016,23,0.898013    ",
  "15042016,23,0.903609    ",
  "16042016,23,0.912827    ",
  "17042016,23,0.927098    ",
  "18042016,23,0.917130    ",
  "19042016,23,0.924094    ",
  "20042016,23,0.951444    ",
  "21042016,23,0.965599    ",
  "22042016,23,0.912480    ",
  "23042016,23,0.895554    ",
  "24042016,23,0.903807    ",
  "25042016,23,0.901850    ",
  "26042016,23,0.912165    ",
  "27042016,23,0.917750    ",
  "28042016,23,0.935242    ",
  "29042016,23,0.951913    ",
  "30042016,23,0.927160    ",
  "01052016,23,0.943811    ",
  "02052016,23,0.897388    ",
  "03052016,23,0.901410    ",
  "04052016,23,0.977341    ",
  "05052016,23,0.930305    ",
  "06052016,23,0.894134    ",
  "07052016,23,0.862451    ",
  "08052016,23,0.905636    ",
  "09052016,23,0.886463    ",
  "10052016,23,0.860881    ",
  "11052016,23,0.868558    ",
  "12052016,23,0.869709    ",
  "13052016,23,0.879589    ",
  "14052016,23,0.884853    ",
  "15052016,23,0.882387    ",
  "16052016,23,0.892936    ",
  "17052016,23,0.825145    ",
  "18052016,23,0.694486    ",
  "19052016,23,0.873818    ",
  "20052016,23,0.878225    ",
  "21052016,23,0.878078    ",
  "22052016,23,0.882108    ",
  "23052016,23,0.882265    ",
  "24052016,23,0.869724    ",
  "25052016,23,0.845536    ",
  "26052016,23,0.869547    ",
  "27052016,23,0.818007    ",
  "28052016,23,0.775234    ",
  "29052016,23,0.884018    ",
  "30052016,23,0.816625    ",
  "31052016,23,0.867032    ",
  "01062016,23,0.874700    ",
  "02062016,23,0.880007    ",
  "03062016,23,0.880426    ",
  "04062016,23,0.885012    ",
  "05062016,23,0.889055    ",
  "06062016,23,0.890951    ",
  "07062016,23,0.859103    ",
  "08062016,23,0.873869    ",
  "09062016,23,0.884626    ",
  "10062016,23,0.896390    ",
  "11062016,23,0.902788    ",
  "12062016,23,0.897016    ",
  "13062016,23,0.897680    ",
  "14062016,23,0.897456    ",
  "15062016,23,0.897302    ",
  "16062016,23,0.898118    ",
  "17062016,23,0.897711    ",
  "18062016,23,0.896380    ",
  "19062016,23,0.847139    ",
  "20062016,23,0.792261    ",
  "21062016,23,0.744220    ",
  "22062016,23,0.641165    ",
  "23062016,23,0.238726    ",
  "24062016,23,0.157712    ",
  "25062016,23,-0.130578   ",
  "26062016,23,-0.161135   ",
  "27062016,23,-0.167744   ",
  "28062016,23,-0.192503   ",
  "29062016,23,-0.189429   ",
  "30062016,23,-0.215659   ",
  "01072016,23,-0.230866   ",
  "02072016,23,-0.249507   ",
  "03072016,23,-0.249565   ",
  "04072016,23,-0.262408   ",
  "05072016,23,-0.270081   ",
  "06072016,23,-0.279906   ",
  "07072016,23,-0.286102   ",
  "08072016,23,-0.292327   ",
  "09072016,23,-0.300834   ",
  "10072016,23,-0.304848   ",
  "11072016,23,-0.314632   ",
  "12072016,23,-0.315711   ",
  "13072016,23,-0.297080   ",
  "14072016,23,-0.285249   ",
  "15072016,23,-0.279831   ",
  "16072016,23,-0.263656   ",
  "17072016,23,-0.246617   ",
  "18072016,23,-0.220854   ",
  "19072016,23,-0.200635   ",
  "20072016,23,-0.185350   ",
  "21072016,23,-0.175160   ",
  "22072016,23,-0.151390   ",
  "23072016,23,-0.134813   ",
  "24072016,23,-0.122510   ",
  "25072016,23,-0.113663   ",
  "26072016,23,-0.108560   ",
  "27072016,23,-0.108251   ",
  "28072016,23,-0.115665   ",
  "29072016,23,-0.124711   ",
  "30072016,23,-0.136648   ",
  "31072016,23,-0.147505   ",
  "01082016,23,-0.149058   ",
  "02082016,23,-0.151780   ",
  "03082016,23,-0.158502   ",
  "04082016,23,-0.167761   ",
  "05082016,23,-0.176287   ",
  "06082016,23,-0.185615   ",
  "07082016,23,-0.190003   ",
  "08082016,23,-0.186368   ",
  "09082016,23,-0.183589   ",
  "10082016,23,-0.173680   ",
  "11082016,23,-0.150381   ",
  "12082016,23,-0.122229   ",
  "13082016,23,-0.089393   ",
  "14082016,23,-0.066207   ",
  "15082016,23,-0.047175   ",
  "16082016,23,-0.027101   ",
  "17082016,23,0.001170    ",
  "18082016,23,0.039912    ",
  "19082016,23,0.106603    ",
  "20082016,23,0.167334    ",
  "21082016,23,0.218204    ",
  "22082016,23,0.260054    ",
  "23082016,23,0.302101    ",
  "24082016,23,0.335605    ",
  "25082016,23,0.376005    ",
  "26082016,23,0.427081    ",
  "27082016,23,0.471664    ",
  "28082016,23,0.511756    ",
  "29082016,23,0.548298    ",
  "30082016,23,0.603619    ",
  "31082016,23,0.640154    ",
  "01092016,23,0.667200    ",
  "02092016,23,0.712057    ",
  "03092016,23,0.730774    ",
  "04092016,23,0.762303    ",
  "05092016,23,0.791664    ",
  "06092016,23,0.816714    ",
  "07092016,23,0.831476    ",
  "08092016,23,0.846911    ",
  "09092016,23,0.869354    ",
  "10092016,23,0.887145    ",
  "11092016,23,0.905861    ",
  "12092016,23,0.898025    ",
  "13092016,23,0.898561    ",
  "14092016,23,0.898507    ",
  "15092016,23,0.898730    ",
  "16092016,23,0.899201    ",
  "17092016,23,0.899420    ",
  "18092016,23,0.899392    ",
  "19092016,23,0.899363    ",
  "20092016,23,0.899363    ",
  "21092016,23,0.898895    ",
  "22092016,23,0.899377    ",
  "23092016,23,0.899381    ",
  "24092016,23,0.899369    ",
  "25092016,23,0.899369    ",
  "26092016,23,0.899372    ",
  "27092016,23,0.899370    ",
  "28092016,23,0.899370    ",
  "29092016,23,0.899379    ",
  "30092016,23,0.899377    ",
  "01102016,23,0.899375    ",
  "02102016,23,0.899377    ",
  "03102016,23,0.899373    ",
  "04102016,23,0.899376    ",
  "05102016,23,0.899378    ",
  "06102016,23,0.899145    ",
  "07102016,23,0.876596    ",
  "08102016,23,0.899082    ",
  "09102016,23,0.899371    ",
  "10102016,23,0.895837    ",
  "11102016,23,0.899358    ",
  "12102016,23,0.896917    ",
  "13102016,23,0.899447    ",
  "14102016,23,0.863238    ",
  "15102016,23,0.873326    ",
  "16102016,23,0.896398    ",
  "17102016,23,0.873132    ",
  "18102016,23,0.894933    ",
  "19102016,23,0.895685    ",
  "20102016,23,0.865714    ",
  "21102016,23,0.882060    ",
  "22102016,23,0.890674    ",
  "23102016,23,0.893399    ",
  "24102016,23,0.813735    ",
  "25102016,23,0.798958    ",
  "26102016,23,0.880389    ",
  "27102016,23,0.741579    ",
  "28102016,23,0.711785    ",
  "29102016,23,0.855402    ",
  "30102016,23,0.854340    ",
  "31102016,23,0.807808    ",
  "01112016,23,0.745079    ",
  "02112016,23,0.812930    ",
  "03112016,23,0.814089    ",
  "04112016,23,0.880723    ",
  "05112016,23,0.798367    ",
  "06112016,23,0.871464    ",
  "07112016,23,0.888897    ",
  "08112016,23,0.869867    ",
  "09112016,23,0.887917    ",
  "10112016,23,0.868678    ",
  "11112016,23,0.864517    ",
  "12112016,23,0.878531    ",
  "13112016,23,0.830401    ",
  "14112016,23,0.726142    ",
  "15112016,23,0.617964    ",
  "16112016,23,0.141111    ",
  "17112016,23,-0.041755   ",
  "18112016,23,-0.107422   ",
  "19112016,23,-0.103700   ",
  "20112016,23,-0.138118   ",
  "21112016,23,-0.164078   ",
  "22112016,23,-0.190549   ",
  "23112016,23,-0.191047   ",
  "24112016,23,-0.187880   ",
  "25112016,23,-0.186013   ",
  "26112016,23,-0.187100   ",
  "27112016,23,-0.190988   ",
  "28112016,23,-0.188752   ",
  "29112016,23,-0.187456   ",
  "30112016,23,-0.186526   ",
  "01122016,23,-0.187001   ",
  "02122016,23,-0.182445   ",
  "03122016,23,-0.179953   ",
  "04122016,23,-0.180305   ",
  "05122016,23,-0.181177   ",
  "06122016,23,-0.184701   ",
  "07122016,23,-0.181579   ",
  "08122016,23,-0.192495   ",
  "09122016,23,-0.204165   ",
  "10122016,23,-0.219398   ",
  "11122016,23,-0.224525   ",
  "12122016,23,-0.217256   ",
  "13122016,23,-0.218930   ",
  "14122016,23,-0.219810   ",
  "15122016,23,-0.216711   ",
  "16122016,23,-0.244493   ",
  "17122016,23,-0.251745   ",
  "18122016,23,-0.246339   ",
  "19122016,23,-0.240272   ",
  "20122016,23,-0.235390   ",
  "21122016,23,-0.233024   ",
  "22122016,23,-0.227190   ",
  "23122016,23,-0.229797   ",
  "24122016,23,-0.234224   ",
  "25122016,23,-0.225309   ",
  "26122016,23,-0.216935   ",
  "27122016,23,-0.210292   ",
  "28122016,23,-0.203410   ",
  "29122016,23,-0.196888   ",
  "30122016,23,-0.192361   ",
  "31122016,23,-0.193337   " ;

 me2016f =
  "31052016  0  0  0  0  1.68124  0  1.68124  0  0  0  0  0  0  0  0  0  0  0  0  0.02  0.76  0  0  1  0  0                        ",
  "16062016  0  0  0  0  0  0  6.72495  0  0  0  0  0  0  0  0  0  0  0  0  0.02  0.76  0  0  1  0  0                              ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                ",
  "                                                                                                                                " ;
}
