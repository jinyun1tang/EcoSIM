netcdf Blodget_pft_20240622.ENF {
dimensions:
	ntopou = 1 ;
	nchar1 = 10 ;
	nchar2 = 10 ;
	ncharmgnt = 128 ;
	maxpfts = 5 ;
	maxpmgt = 24 ;
	year = UNLIMITED ; // (2 currently)
variables:
	int NH1(ntopou) ;
		NH1:long_name = "Starting column from the west for a topo unit" ;
		NH1:units = "None" ;
	int NV1(ntopou) ;
		NV1:long_name = "Ending column at the east for a topo unit" ;
		NV1:units = "None" ;
	int NH2(ntopou) ;
		NH2:long_name = "Starting row from the north  for a topo unit" ;
		NH2:units = "None" ;
	int NV2(ntopou) ;
		NV2:long_name = "Ending row at the south  for a topo unit" ;
		NV2:units = "None" ;
	int NZ(ntopou) ;
		NZ:long_name = "Number of pfts on a topo unit" ;
		NZ:units = "None" ;
	short nmgnts(year, ntopou, maxpfts) ;
		nmgnts:long_name = "Number of managements for a given pft in in given topo unit in a year" ;
	char pft_type(year, ntopou, maxpfts, nchar1) ;
	char pft_pltinfo(year, ntopou, maxpfts, ncharmgnt) ;
		pft_pltinfo:long_name = "string containing planting information" ;
	char pft_mgmt(year, ntopou, maxpfts, maxpmgt, ncharmgnt) ;
		pft_mgmt:long_name = "string containing plant management information" ;
	int pft_dflag ;
		pft_dflag:long_name = "Flag for plant management data" ;
		pft_dflag:flags = "-1 no pft data, 0 only plantation information, 1 transient pft data" ;

// global attributes:
		:description = "PFT input data created on 2024/06/22/11:44:43\n",
			" use READ(tline,*)DY,PPI(NZ,NY,NX),SDPTHI(NZ,NY,NX) to read planting information from pft_pltinfo; use READ(tline,*)DY,ICUT,JCUT,HCUT,PCUT,ECUT11,ECUT12,ECUT13,ECUT14,ECUT21,ECUT22,ECUT23,ECUT24 to read management information from pft_mgmt" ;
data:

 NH1 = 1 ;

 NV1 = 1 ;

 NH2 = 1 ;

 NV2 = 1 ;

 NZ = 2 ;

 nmgnts =
  0, 0, _, _, _,
  12, 12, _, _, _ ;

 pft_type =
  "ndlf34",
  "dfir34",
  "",
  "",
  "",
  "ndlf34",
  "dfir34",
  "",
  "",
  "" ;

 pft_pltinfo =
  "01019999 0.015 0.011                                                                                                            ",
  "01019999 0.015 0.011                                                                                                            ",  
  "",
  "",
  "",
  "01010000 0.015 0.011                                                                                                            ",
  "01010000 0.015 0.011                                                                                                            ",  
  "",
  "",
  "" ;

 pft_mgmt =
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "31010000 0 0 1000 0.00083 1 1 1 0 0 0 0 0                                                                                       ",
  "28020000 0 0 1000 0.00083 1 1 1 0 0 0 0 0                                                                                       ",
  "31030000 0 0 1000 0.00083 1 1 1 0 0 0 0 0                                                                                       ",
  "30040000 0 0 1000 0.00083 1 1 1 0 0 0 0 0                                                                                       ",
  "31050000 0 0 1000 0.00083 1 1 1 0 0 0 0 0                                                                                       ",
  "30060000 0 0 1000 0.00083 1 1 1 0 0 0 0 0                                                                                       ",
  "31070000 0 0 1000 0.00083 1 1 1 0 0 0 0 0                                                                                       ",
  "31080000 0 0 1000 0.00083 1 1 1 0 0 0 0 0                                                                                       ",
  "30090000 0 0 1000 0.00083 1 1 1 0 0 0 0 0                                                                                       ",
  "31100000 0 0 1000 0.00083 1 1 1 0 0 0 0 0                                                                                       ",
  "30110000 0 0 1000 0.00083 1 1 1 0 0 0 0 0                                                                                       ",
  "30120000 0 0 1000 0.00083 1 1 1 0 0 0 0 0                                                                                       ",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "31010000 0 0 1000 0.00083 1 1 1 0 0 0 0 0                                                                                       ",
  "28020000 0 0 1000 0.00083 1 1 1 0 0 0 0 0                                                                                       ",
  "31030000 0 0 1000 0.00083 1 1 1 0 0 0 0 0                                                                                       ",
  "30040000 0 0 1000 0.00083 1 1 1 0 0 0 0 0                                                                                       ",
  "31050000 0 0 1000 0.00083 1 1 1 0 0 0 0 0                                                                                       ",
  "30060000 0 0 1000 0.00083 1 1 1 0 0 0 0 0                                                                                       ",
  "31070000 0 0 1000 0.00083 1 1 1 0 0 0 0 0                                                                                       ",
  "31080000 0 0 1000 0.00083 1 1 1 0 0 0 0 0                                                                                       ",
  "30090000 0 0 1000 0.00083 1 1 1 0 0 0 0 0                                                                                       ",
  "31100000 0 0 1000 0.00083 1 1 1 0 0 0 0 0                                                                                       ",
  "30110000 0 0 1000 0.00083 1 1 1 0 0 0 0 0                                                                                       ",
  "30120000 0 0 1000 0.00083 1 1 1 0 0 0 0 0                                                                                       ",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "" ;

 pft_dflag = 0 ;
}
